* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

* Placeholder for "condiode", which probably represents the parasitic
* well-to-substrate diode, although it does not take any parameters.
.SUBCKT sky130_fd_io__condiode NEG POS
.ENDS

.SUBCKT sky130_fd_io__gnd2gnd_120x2_lv_isosub BDY2_B2B SRC_BDY_LVC1 VSSD
D0 SRC_BDY_LVC1 BDY2_B2B sky130_fd_pr__diode_pd2nw_05v5 area=90E+12 pj=132E+6
D1 BDY2_B2B SRC_BDY_LVC1 sky130_fd_pr__diode_pd2nw_05v5 area=90E+12 pj=132E+6
.ENDS

.SUBCKT sky130_fd_io__amuxsplitv2_delay ENABLE_VDDA_H HLD_VDDA_H_N HOLD RESET
+ VCC_IO VGND
*.PININFO ENABLE_VDDA_H:I HLD_VDDA_H_N:I HOLD:O RESET:O VCC_IO:B
*.PININFO VGND:B
XI33 enable_vdda_switch hld_vdda_h_n_switch RESET VGND VCC_IO
+ sky130_fd_io__hvsbt_nand2
XI29 hld_vdda_h_n_switch hld_vdda_h VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5
+ m=2 w=3.0 l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI28 hld_vdda_h HLD_VDDA_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=3.0 l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI12 enable_vdda_switch enable_vdda_h_n VCC_IO VCC_IO
+ sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
XI13 enable_vdda_h_n ENABLE_VDDA_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5
+ m=1 w=3.0 l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI36 HOLD RESET VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI31 hld_vdda_h_n_switch hld_vdda_h VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=2
+ w=1.0 l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI30 hld_vdda_h HLD_VDDA_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI14 enable_vdda_switch enable_vdda_h_n VGND VGND sky130_fd_pr__nfet_g5v0d10v5
+ m=2 w=1.0 l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI15 enable_vdda_h_n ENABLE_VDDA_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=1.0 l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI37 HOLD RESET VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__amuxsplitv2_delay

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__amuxsplitv2_switch AMUXBUS_L AMUXBUS_R NGATE_SL_H
+ NGATE_SR_H NMID_H PGATE_SL_H_N PGATE_SR_H_N VDDA VSSA
*.PININFO AMUXBUS_L:B AMUXBUS_R:B NGATE_SL_H:I NGATE_SR_H:I NMID_H:I
*.PININFO PGATE_SL_H_N:I PGATE_SR_H_N:I VDDA:B VSSA:B
xI20 mid VDDA sky130_fd_io__condiode
xI19 VSSA VDDA sky130_fd_io__condiode
XI18 VSSA nmid_h_s sky130_fd_io__res75only_small
XI1 AMUXBUS_L NGATE_SL_H mid mid sky130_fd_pr__nfet_g5v0d10v5 m=30 w=10.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 mid NGATE_SR_H AMUXBUS_R mid sky130_fd_pr__nfet_g5v0d10v5 m=30 w=10.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI4 mid NMID_H nmid_h_s VSSA sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI0 mid PGATE_SL_H_N AMUXBUS_L VDDA sky130_fd_pr__pfet_g5v0d10v5 m=14 w=10.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI3 AMUXBUS_R PGATE_SR_H_N mid VDDA sky130_fd_pr__pfet_g5v0d10v5 m=14 w=10.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__amuxsplitv2_switch

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__amuxsplitv2_switch_levelshifter FBK FBK_N HOLD RESET
+ SWITCH_LV SWITCH_LV_N VGND VPWR_HV VPWR_LV
*.PININFO FBK:O FBK_N:O HOLD:I RESET:I SWITCH_LV:I SWITCH_LV_N:I
*.PININFO VGND:B VPWR_HV:B VPWR_LV:B
XI184 FBK RESET VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI183 net97 VPWR_LV net109 VGND sky130_fd_pr__nfet_05v0_nvt m=4 w=1.0 l=0.9
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI18 FBK HOLD net105 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI182 net105 VPWR_LV net117 VGND sky130_fd_pr__nfet_05v0_nvt m=4 w=1.0 l=0.9
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI16 net109 SWITCH_LV VGND VGND sky130_fd_pr__nfet_01v8_lvt m=4 w=1.0 l=0.15
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI15 FBK_N HOLD net97 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI19 net117 SWITCH_LV_N VGND VGND sky130_fd_pr__nfet_01v8_lvt m=4 w=1.0 l=0.15
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI185 FBK_N FBK VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI20 FBK FBK_N VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__amuxsplitv2_switch_levelshifter

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__amuxsplitv2_switch_s0 HOLD IN_LV OUT_H RESET VCCD VDDA
+ VSSA VSSD
*.PININFO HOLD:I IN_LV:I OUT_H:O RESET:I VCCD:B VDDA:B VSSA:B VSSD:B
XI0 net17 net13 HOLD RESET in_lv_i in_lv_n VSSA VDDA VCCD
+ sky130_fd_io__amuxsplitv2_switch_levelshifter
XI22 in_lv_n IN_LV VSSD VSSD sky130_fd_pr__nfet_01v8 m=1 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI21 in_lv_i in_lv_n VSSD VSSD sky130_fd_pr__nfet_01v8 m=1 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI16 OUT_H net13 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI20 in_lv_n IN_LV VCCD VCCD sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI19 in_lv_i in_lv_n VCCD VCCD sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI15 OUT_H net13 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__amuxsplitv2_switch_s0

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__amuxsplitv2_switch_sl HOLD IN_LV OUT_H OUT_H_N RESET VCCD
+ VDDA VSSA VSSD VSWITCH
*.PININFO HOLD:I IN_LV:I OUT_H:O OUT_H_N:O RESET:I VCCD:B VDDA:B
*.PININFO VSSA:B VSSD:B VSWITCH:B
XI0 net39 net35 HOLD RESET in_lv_i in_lv_n VSSA VDDA VCCD
+ sky130_fd_io__amuxsplitv2_switch_levelshifter
XI1 net48 net44 HOLD RESET in_lv_i in_lv_n VSSA VSWITCH VCCD
+ sky130_fd_io__amuxsplitv2_switch_levelshifter
XI14 OUT_H net44 VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI15 OUT_H_N net39 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI19 in_lv_i in_lv_n VCCD VCCD sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI20 in_lv_n IN_LV VCCD VCCD sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI13 OUT_H net44 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI16 OUT_H_N net39 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI21 in_lv_i in_lv_n VSSD VSSD sky130_fd_pr__nfet_01v8 m=1 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI22 in_lv_n IN_LV VSSD VSSD sky130_fd_pr__nfet_01v8 m=1 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__amuxsplitv2_switch_sl

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__amx_inv1 A Y VDA VSSA
*.PININFO A:I Y:O VDA:I VSSA:I
XI92 Y A VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI54 Y A VDA VDA sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__amx_inv1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_cclat DRVHI_H DRVLO_H_N OE_H_N PD_DIS_H PU_DIS_H
+ VCC_IO VGND
*.PININFO DRVHI_H:O DRVLO_H_N:O OE_H_N:I PD_DIS_H:I PU_DIS_H:I
*.PININFO VCC_IO:I VGND:I
Xnor3_q0 oe_i_h_n DRVHI_H PD_DIS_H n1 VCC_IO VGND VGND
+ sky130_fd_io__com_cclat_hvnor3
Xnand3_q0 oe_i_h DRVLO_H_N pu_dis_h_n n0 VCC_IO VGND VGND
+ sky130_fd_io__com_cclat_hvnand3
Xinv_oe1_q0 OE_H_N oe_i_h VCC_IO VGND VGND sky130_fd_io__com_cclat_inv_in
Xinv_oe2_q0 oe_i_h oe_i_h_n VCC_IO VGND VGND sky130_fd_io__com_cclat_inv_in
Xinv_pudis_q0 PU_DIS_H pu_dis_h_n VCC_IO VGND VGND
+ sky130_fd_io__com_cclat_inv_in
Xinv_out_q0 n1 DRVLO_H_N VCC_IO VGND VGND sky130_fd_io__com_cclat_inv_out
Xinv_out_1_q0 n0 DRVHI_H VCC_IO VGND VGND sky130_fd_io__com_cclat_inv_out
.ENDS sky130_fd_io__com_cclat

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_cclat_hvnand3 IN0 IN1 IN2 OUT VCC_IO VGND VNB
*.PININFO IN0:I IN1:I IN2:I OUT:O VCC_IO:I VGND:I VNB:I
Xmp0_q0 OUT IN0 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmp2_q0 OUT IN2 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmp1_q0 OUT IN1 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmn2_q0 OUT IN2 n1 VNB sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmn0_q0 n0 IN0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=4 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmn1_q0 n1 IN1 n0 VNB sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_cclat_hvnand3

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_cclat_hvnor3 IN0 IN1 IN2 OUT VCC_IO VGND VNB
*.PININFO IN0:I IN1:I IN2:I OUT:O VCC_IO:I VGND:I VNB:I
Xmp0_q0 n<0> IN0 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=8 w=5.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmp2_q0 OUT IN2 n<1> VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmp1_q0 n<1> IN1 n<0> VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmn0_q0 OUT IN0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmn2_q0 OUT IN2 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmn1_q0 OUT IN1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_cclat_hvnor3

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_cclat_i2c_fix DRVHI_H DRVLO_H_N OE_H PD_DIS_H PU_DIS_H
+ VCC_IO VGND
*.PININFO DRVHI_H:O DRVLO_H_N:O OE_H:I PD_DIS_H:I PU_DIS_H:I VCC_IO:I
*.PININFO VGND:I
Xnor3_q0 oe_i_h_n DRVHI_H PD_DIS_H n1 VCC_IO VGND VGND
+ sky130_fd_io__com_cclat_hvnor3
Xnand3_q0 OE_H DRVLO_H_N pu_dis_h_n n0 VCC_IO VGND VGND
+ sky130_fd_io__com_cclat_hvnand3
Xinv_oe2_q0 OE_H oe_i_h_n VCC_IO VGND VGND sky130_fd_io__com_cclat_inv_in
Xinv_pudis_q0 PU_DIS_H pu_dis_h_n VCC_IO VGND VGND
+ sky130_fd_io__com_cclat_inv_in
Xinv_out_q0 n1 DRVLO_H_N VCC_IO VGND VGND sky130_fd_io__com_cclat_inv_out
Xinv_out_1_q0 n0 DRVHI_H VCC_IO VGND VGND sky130_fd_io__com_cclat_inv_out
.ENDS sky130_fd_io__com_cclat_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_cclat_inv_in IN OUT VCC_IO VGND VNB
*.PININFO IN:I OUT:O VCC_IO:I VGND:I VNB:I
Xmp1_q0 OUT IN VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmn1_q0 OUT IN VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_cclat_inv_in

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_cclat_inv_out IN OUT VCC_IO VGND VNB
*.PININFO IN:I OUT:O VCC_IO:I VGND:I VNB:I
XI1 OUT IN VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=6 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 OUT IN VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=6 w=3.0 l=0.6 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_cclat_inv_out

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_ctl_ls HLD_H_N IN OUT_H OUT_H_N RST_H SET_H VCC_IO
+ VGND VPWR
*.PININFO HLD_H_N:I IN:I OUT_H:O OUT_H_N:O RST_H:I SET_H:I VCC_IO:I
*.PININFO VGND:I VPWR:I
XI14 OUT_H_N fbk VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI34 in_i in_i_n VPWR VPWR sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI29 in_i_n IN VPWR VPWR sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI11 OUT_H fbk_n VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 fbk fbk_n VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 fbk_n fbk VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI13 OUT_H_N fbk VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmnset_q0 fbk_n SET_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI32 in_i in_i_n VGND VGND sky130_fd_pr__nfet_01v8 m=1 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 OUT_H fbk_n VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI58 net130 VPWR net94 VGND sky130_fd_pr__nfet_05v0_nvt m=4 w=1.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmnrst_q0 fbk RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI59 net122 VPWR net98 VGND sky130_fd_pr__nfet_05v0_nvt m=4 w=1.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 fbk_n HLD_H_N net122 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI27 in_i_n IN VGND VGND sky130_fd_pr__nfet_01v8 m=1 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI5 fbk HLD_H_N net130 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI4 fbk_n fbk VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI3 fbk fbk_n VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.75 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI8 net98 in_i VGND VGND sky130_fd_pr__nfet_01v8_lvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI7 net94 in_i_n VGND VGND sky130_fd_pr__nfet_01v8_lvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_ctl_ls

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_inv_x1_dnw IN OUT VGND VPWR
*.PININFO IN:I OUT:O VGND:I VPWR:I
XI1 OUT IN VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 OUT IN VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_inv_x1_dnw

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_nand2_dnw IN0 IN1 OUT VGND VPWR
*.PININFO IN0:I IN1:I OUT:O VGND:I VPWR:I
XI3 OUT IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI5 OUT IN1 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN1 net25 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 net25 IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_nand2_dnw

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_nor2_dnw IN0 IN1 OUT VGND VPWR
*.PININFO IN0:I IN1:I OUT:O VGND:I VPWR:I
XI3 net17 IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 OUT IN1 net17 VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 OUT IN1 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_nor2_dnw

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_pad PAD VGND_IO
*.PININFO PAD:B VGND_IO:B
.ENDS sky130_fd_io__com_pad

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_pddrvr_unit_2_5 ND NGIN NS
*.PININFO ND:B NGIN:I NS:B
Xndrv_q0 ND NGIN NS NS sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_pddrvr_unit_2_5

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_pdpredrvr_pbias DRVLO_H_N EN_H EN_H_N PBIAS PD_H
+ PDEN_H_N VCC_IO VGND_IO
*.PININFO DRVLO_H_N:I EN_H:I EN_H_N:I PBIAS:O PD_H:I PDEN_H_N:I
*.PININFO VCC_IO:I VGND_IO:I
XI27 n<0> PD_H EN_H_N sky130_fd_io__tk_opto
XE1 n<1> n<0> sky130_fd_io__tk_em1o
XE2 PBIAS pbias1 sky130_fd_io__tk_em1o
XE3 pbias1 net88 sky130_fd_io__tk_em1s
XE4 net108 PBIAS sky130_fd_io__tk_em1s
XE6 PBIAS net84 sky130_fd_io__tk_em1s
XE5 n<101> bias_g sky130_fd_io__tk_em1s
XI47 PBIAS bias_g VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.0 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI24 n<1> DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI18 bias_g DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI23 n<0> n<0> n<1> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI13 drvlo_i_h DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI20 bias_g n<1> VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI19 bias_g EN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI34 net157 bias_g VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI36 net108 bias_g VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.0 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI38 n<1> PDEN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI48 n<100> PD_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=4.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI41 n<101> PD_H n<100> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=4.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI44 PBIAS PBIAS pbias1 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=8 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI45 pbias1 pbias1 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=8 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI15 net183 EN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI16 net171 n<0> net183 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 PBIAS EN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 drvlo_i_h DRVLO_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI17 bias_g DRVLO_H_N net171 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI14 PBIAS drvlo_i_h VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI33 N0 VGND_IO VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=8.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI32 net161 net161 N0 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI31 net157 net157 net161 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI30 net88 N0 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=8 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI43 net84 bias_g VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=4.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI40 N0 drvlo_i_h VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_pdpredrvr_pbias

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_pdpredrvr_strong_slow DRVLO_H_N PD_H PDEN_H_N VCC_IO
+ VGND_IO
*.PININFO DRVLO_H_N:I PD_H:O PDEN_H_N:I VCC_IO:I VGND_IO:I
XI26 PD_H PDEN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI25 PD_H DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI24 net25 PDEN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI23 PD_H DRVLO_H_N net25 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_pdpredrvr_strong_slow

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_pdpredrvr_weak DRVLO_H_N PD_H PDEN_H_N VCC_IO VGND_IO
*.PININFO DRVLO_H_N:I PD_H:O PDEN_H_N:I VCC_IO:I VGND_IO:I
XI26 PD_H PDEN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI25 PD_H DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI24 net25 PDEN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI23 PD_H DRVLO_H_N net25 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_pdpredrvr_weak

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_pudrvr_strong_slow PAD PU_H_N VCC_IO VGND_IO VPB_DRVR
*.PININFO PAD:O PU_H_N:I VCC_IO:I VGND_IO:I VPB_DRVR:I
Xpdrv_q0 PAD PU_H_N VCC_IO VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=8 w=7.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_pudrvr_strong_slow

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_pudrvr_weak PAD PU_H_N VCC_IO VGND_IO VPB_DRVR
*.PININFO PAD:O PU_H_N:I VCC_IO:I VGND_IO:I VPB_DRVR:I
Xpdrv_q0 PAD PU_H_N VCC_IO VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=4 w=7.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI29 PAD PU_H_N VCC_IO VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_pudrvr_weak

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_pupredrvr_nbias DRVHI_H EN_H EN_H_N NBIAS PU_H_N
+ PUEN_H VCC_IO VGND_IO
*.PININFO DRVHI_H:I EN_H:I EN_H_N:I NBIAS:O PU_H_N:I PUEN_H:I VCC_IO:I
*.PININFO VGND_IO:I
XI36 n<2> PU_H_N EN_H sky130_fd_io__tk_opto
XE5 NBIAS net88 sky130_fd_io__tk_em1s
XE4 n<6> net153 sky130_fd_io__tk_em1s
XE7 bias_g net90 sky130_fd_io__tk_em1s
XE6 net141 NBIAS sky130_fd_io__tk_em1s
XE1 n<2> n<1> sky130_fd_io__tk_em1o
XE2 n<6> NBIAS sky130_fd_io__tk_em1o
XI34 n<1> DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI32 n<1> n<2> n<2> VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI31 bias_g n<1> VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=4 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI30 bias_g DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI29 bias_g EN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI21 NBIAS bias_g VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.0 l=0.8
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 drvhi_i_h_n DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI47 n<7> bias_g VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI49 net88 bias_g VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.0 l=0.8
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI50 n<1> PUEN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI56 VCC_IO PU_H_N net90 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=8.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI19 n<6> n<6> VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=4 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI20 NBIAS NBIAS n<6> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=4 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI28 bias_g DRVHI_H n<3> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI27 n<3> n<2> n<4> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI26 n<4> EN_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI13 drvhi_i_h_n DRVHI_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI24 NBIAS EN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI53 vccio_2vtn drvhi_i_h_n VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=3.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI25 NBIAS drvhi_i_h_n VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI40 vccio_2vtn VCC_IO VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI39 net153 vccio_2vtn VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=4 w=3.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI44 n<8> n<8> vccio_2vtn VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI41 n<7> n<7> n<8> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI54 net141 bias_g VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=4.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_pupredrvr_nbias

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_pupredrvr_strong_slow DRVHI_H PU_H_N PUEN_H VCC_IO
+ VGND_IO
*.PININFO DRVHI_H:I PU_H_N:O PUEN_H:I VCC_IO:I VGND_IO:I
XI3 PU_H_N DRVHI_H net17 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI39 net17 PUEN_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI38 PU_H_N PUEN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI37 PU_H_N DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=3 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_pupredrvr_strong_slow

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_pupredrvr_weak DRVHI_H PU_H_N PUEN_H VCC_IO VGND_IO
*.PININFO DRVHI_H:I PU_H_N:O PUEN_H:I VCC_IO:I VGND_IO:I
XI3 PU_H_N DRVHI_H net21 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI39 net21 PUEN_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI38 PU_H_N PUEN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI37 PU_H_N DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__com_pupredrvr_weak

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_res_strong_slow RA RB VGND_IO
*.PININFO RA:B RB:B VGND_IO:I
XI28 net34 net30 sky130_fd_io__tk_em1s
RI32 RB net30 sky130_fd_pr__res_generic_po W=2 L=2 m=1
RI29 net30 net34 sky130_fd_pr__res_generic_po W=2 L=3 m=1
Rr1 net34 RA sky130_fd_pr__res_generic_po W=2 L=5 m=1
.ENDS sky130_fd_io__com_res_strong_slow

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_res_weak RA RB VGND_IO
*.PININFO RA:B RB:B VGND_IO:I
Xe9_q0 n<0> n<1> sky130_fd_io__tk_em1s
Xe11_q0 n<2> n<3> sky130_fd_io__tk_em1s
Xe10_q0 n<1> n<2> sky130_fd_io__tk_em1s
Xe12_q0 n<3> RB sky130_fd_io__tk_em1s
Xe13_q0 n<4> n<0> sky130_fd_io__tk_em1s
Xe14_q0 n<5> n<4> sky130_fd_io__tk_em1o
RI84 n<0> n<1> sky130_fd_pr__res_generic_po W=0.8 L=1.5 m=1
RI62 n<3> RB sky130_fd_pr__res_generic_po W=0.8 L=1.5 m=1
RI82 n<2> n<3> sky130_fd_pr__res_generic_po W=0.8 L=1.5 m=1
RI85 RA net64 sky130_fd_pr__res_generic_po W=0.8 L=50 m=1
RI83 n<1> n<2> sky130_fd_pr__res_generic_po W=0.8 L=1.5 m=1
RI116 net64 n<5> sky130_fd_pr__res_generic_po W=0.8 L=12 m=1
RI104 n<4> n<0> sky130_fd_pr__res_generic_po W=0.8 L=6 m=1
RI134 n<5> n<4> sky130_fd_pr__res_generic_po W=0.8 L=6 m=1
.ENDS sky130_fd_io__com_res_weak

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__com_xres_weak_pu RA RB VGND_IO
*.PININFO RA:B RB:B VGND_IO:I
Xe9_q0 n<0> n<1> sky130_fd_io__tk_em1s
Xe11_q0 n<2> n<3> sky130_fd_io__tk_em1s
Xe10_q0 n<1> n<2> sky130_fd_io__tk_em1s
Xe12_q0 n<3> RB sky130_fd_io__tk_em1s
Xe13_q0 n<4> n<0> sky130_fd_io__tk_em1s
Xe14_q0 n<5> n<4> sky130_fd_io__tk_em1o
RI84 n<0> n<1> sky130_fd_pr__res_generic_po W=0.8 L=1.5 m=1
RI62 n<3> RB sky130_fd_pr__res_generic_po W=0.8 L=1.5 m=1
RI82 n<2> n<3> sky130_fd_pr__res_generic_po W=0.8 L=1.5 m=1
RI85 RA net64 sky130_fd_pr__res_generic_po W=0.8 L=50 m=1
RI83 n<1> n<2> sky130_fd_pr__res_generic_po W=0.8 L=1.5 m=1
RI116 net64 n<5> sky130_fd_pr__res_generic_po W=0.8 L=12 m=1
RI104 n<4> n<0> sky130_fd_pr__res_generic_po W=0.8 L=6 m=1
RI134 n<5> n<4> sky130_fd_pr__res_generic_po W=0.8 L=6 m=1
.ENDS sky130_fd_io__com_xres_weak_pu

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__enh_nand2_1 IN0 IN1 OUT VGND VPWR
*.PININFO IN0:I IN1:I OUT:O VGND:I VPWR:I
XI3 OUT IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=3 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI5 OUT IN1 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=3 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN1 net25 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 net25 IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__enh_nand2_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__enh_nand2_1_sp IN0 IN1 OUT VGND VPWR
*.PININFO IN0:I IN1:I OUT:O VGND:I VPWR:I
XI3 OUT IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI5 OUT IN1 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN1 net25 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 net25 IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__enh_nand2_1_sp

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__enh_nor2_x1 IN0 IN1 OUT VGND VPWR
*.PININFO IN0:I IN1:I OUT:O VGND:I VPWR:I
XI3 net16 IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=2
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 OUT IN1 net16 VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=2
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 OUT IN1 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__enh_nor2_x1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

* Modified by Tim:  The local_5term cells have resistors that overlap, and the resistor
* end terminals must be added to the netlist to make it correct.

.SUBCKT sky130_fd_io__gpio_buf_localesd IN_H OUT_H OUT_VT VCC_IO VGND
+ VTRIP_SEL_H
*.PININFO IN_H:I OUT_H:O OUT_VT:O VCC_IO:B VGND:B VTRIP_SEL_H:I
Xesd_res_q0 IN_H OUT_H sky130_fd_io__res250only_small
Xggnfet2_q0 VGND OUT_VT VGND VCC_IO VGND VCC_IO
+ sky130_fd_io__signal_5_sym_hv_local_5term
Xggnfet6_q0 VGND VCC_IO VGND VCC_IO OUT_H VCC_IO
+ sky130_fd_io__signal_5_sym_hv_local_5term
Xggnfet5_q0 VGND VCC_IO VGND VCC_IO OUT_VT VCC_IO
+ sky130_fd_io__signal_5_sym_hv_local_5term
Xggnfet1_q0 VGND OUT_H VGND VCC_IO VGND VCC_IO
+ sky130_fd_io__signal_5_sym_hv_local_5term
Xhv_passgate_q0 OUT_H VTRIP_SEL_H OUT_VT VGND sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=3.0 l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
.ENDS sky130_fd_io__gpio_buf_localesd

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ctlv2_i2c_fix DM[2] DM[1] DM[0] DM_H[2] DM_H[1]
+ DM_H[0] DM_H_N[2] DM_H_N[1] DM_H_N[0] ENABLE_H ENABLE_INP_H HLD_H_N HLD_I_H_N
+ HLD_I_OVR_H HLD_OVR HYST_TRIM HYST_TRIM_H HYST_TRIM_H_N IB_MODE_SEL[1]
+ IB_MODE_SEL[0] IB_MODE_SEL_H[1] IB_MODE_SEL_H[0] IB_MODE_SEL_H_N[1]
+ IB_MODE_SEL_H_N[0] INP_DIS INP_DIS_H_N OD_I_H_N SLEW_CTL[1] SLEW_CTL[0]
+ SLEW_CTL_H[1] SLEW_CTL_H[0] SLEW_CTL_H_N[1] SLEW_CTL_H_N[0] VCCD VDDIO_Q VSSD
+ VTRIP_SEL VTRIP_SEL_H
*.PININFO DM[2]:I DM[1]:I DM[0]:I DM_H[2]:O DM_H[1]:O DM_H[0]:O
*.PININFO DM_H_N[2]:O DM_H_N[1]:O DM_H_N[0]:O ENABLE_H:I
*.PININFO ENABLE_INP_H:I HLD_H_N:I HLD_I_H_N:O HLD_I_OVR_H:O HLD_OVR:I
*.PININFO HYST_TRIM:I HYST_TRIM_H:O HYST_TRIM_H_N:O IB_MODE_SEL[1]:I
*.PININFO IB_MODE_SEL[0]:I IB_MODE_SEL_H[1]:O IB_MODE_SEL_H[0]:O
*.PININFO IB_MODE_SEL_H_N[1]:O IB_MODE_SEL_H_N[0]:O INP_DIS:I
*.PININFO INP_DIS_H_N:O OD_I_H_N:O SLEW_CTL[1]:I SLEW_CTL[0]:I
*.PININFO SLEW_CTL_H[1]:O SLEW_CTL_H[0]:O SLEW_CTL_H_N[1]:O
*.PININFO SLEW_CTL_H_N[0]:O VCCD:I VDDIO_Q:I VSSD:I VTRIP_SEL:I
*.PININFO VTRIP_SEL_H:O
Xls_bank_q0 DM[2] DM[1] DM[0] DM_H[2] DM_H[1] DM_H[0] DM_H_N[2] DM_H_N[1]
+ DM_H_N[0] HLD_I_H_N HYST_TRIM HYST_TRIM_H HYST_TRIM_H_N IB_MODE_SEL[1]
+ IB_MODE_SEL[0] IB_MODE_SEL_H[1] IB_MODE_SEL_H[0] IB_MODE_SEL_H_N[1]
+ IB_MODE_SEL_H_N[0] INP_DIS net83 INP_DIS_H_N OD_I_H_N SLEW_CTL[1] SLEW_CTL[0]
+ SLEW_CTL_H[1] SLEW_CTL_H[0] SLEW_CTL_H_N[1] SLEW_CTL_H_N[0] startup_rst_h
+ inp_startup_en_h VDDIO_Q VSSD VCCD VTRIP_SEL VTRIP_SEL_H net77
+ sky130_fd_io__gpio_ovtv2_ctl_lsbank_i2c_fix
Xhld_dis_blk_q0 ENABLE_H HLD_H_N HLD_I_H_N HLD_I_OVR_H HLD_OVR OD_I_H_N VDDIO_Q
+ VSSD VCCD sky130_fd_io__gpio_ovtv2_ctl_hld_i2c_fix
XI75 ENABLE_INP_H ENABLE_H startup_rst_h VSSD VDDIO_Q sky130_fd_io__hvsbt_nor
XI56 net109 ENABLE_INP_H net108 VSSD VDDIO_Q sky130_fd_io__hvsbt_nand2
XI77 OD_I_H_N net109 VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
XI57 net108 inp_startup_en_h VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
.ENDS sky130_fd_io__gpio_ctlv2_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_dat_ls HLD_H_N IN OUT_H OUT_H_N RST_H SET_H VCC_IO
+ VGND VPWR_KA
*.PININFO HLD_H_N:I IN:I OUT_H:O OUT_H_N:O RST_H:I SET_H:I VCC_IO:I
*.PININFO VGND:I VPWR_KA:I
XI3 fbk fbk_n VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI4 fbk_n fbk VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI5 fbk HLD_H_N net79 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 fbk_n HLD_H_N net83 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI7 net107 in_i_n VGND VGND sky130_fd_pr__nfet_01v8_lvt m=8 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI8 net103 in_i VGND VGND sky130_fd_pr__nfet_01v8_lvt m=8 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 OUT_H fbk_n VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI13 OUT_H_N fbk VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmnset_q0 fbk_n SET_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmnrst_q0 fbk RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI34 in_i_n IN VGND VGND sky130_fd_pr__nfet_01v8 m=2 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI35 in_i in_i_n VGND VGND sky130_fd_pr__nfet_01v8 m=2 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI31 net83 VPWR_KA net103 VGND sky130_fd_pr__nfet_05v0_nvt m=8 w=1.0 l=0.9
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI30 net79 VPWR_KA net107 VGND sky130_fd_pr__nfet_05v0_nvt m=8 w=1.0 l=0.9
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 fbk_n fbk VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 fbk fbk_n VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI33 in_i in_i_n VPWR_KA VPWR_KA sky130_fd_pr__pfet_01v8_hvt m=1 w=3.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI11 OUT_H fbk_n VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI14 OUT_H_N fbk VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI32 in_i_n IN VPWR_KA VPWR_KA sky130_fd_pr__pfet_01v8_hvt m=1 w=3.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_dat_ls

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_dat_ls_i2c_fix HLD_H_N IN OUT_H_N SET_H SET_H_N
+ VCC_IO VGND VPWR_KA
*.PININFO HLD_H_N:I IN:I OUT_H_N:O SET_H:I SET_H_N:I VCC_IO:I VGND:I
*.PININFO VPWR_KA:I
XI3 fbk fbk_n VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI4 fbk_n fbk VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI5 fbk HLD_H_N net76 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 fbk_n HLD_H_N net80 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI7 net100 in_i_n VGND VGND sky130_fd_pr__nfet_01v8_lvt m=8 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI8 net96 in_i VGND VGND sky130_fd_pr__nfet_01v8_lvt m=8 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI13 OUT_H_N fbk VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmnset_q0 fbk_n SET_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=4 w=0.7 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI34 in_i_n IN VGND VGND sky130_fd_pr__nfet_01v8 m=2 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI35 in_i in_i_n VGND VGND sky130_fd_pr__nfet_01v8 m=2 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI31 net80 VPWR_KA net96 VGND sky130_fd_pr__nfet_05v0_nvt m=8 w=1.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI30 net76 VPWR_KA net100 VGND sky130_fd_pr__nfet_05v0_nvt m=8 w=1.0 l=0.9
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 fbk_n fbk VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 fbk fbk_n VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI33 in_i in_i_n VPWR_KA VPWR_KA sky130_fd_pr__pfet_01v8_hvt m=1 w=3.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI14 OUT_H_N fbk VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI36 fbk SET_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=3 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI32 in_i_n IN VPWR_KA VPWR_KA sky130_fd_pr__pfet_01v8_hvt m=1 w=3.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_dat_ls_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_amux_i2c_fix AMUXBUS_A AMUXBUS_B ANALOG_EN
+ ANALOG_POL ANALOG_SEL ENABLE_VDDA_H ENABLE_VSWITCH_H HLD_I_H_N NGA_PAD_VPMP_H
+ NGB_PAD_VPMP_H NGHS_H OUT PAD PD_CSD_H PGHS_H PU_CSD_H PUG_H[1] PUG_H[0] VCCD
+ VDDA VDDIO VDDIO_Q VPB_DRVR VSSA VSSD VSSIO VSWITCH
*.PININFO AMUXBUS_A:B AMUXBUS_B:B ANALOG_EN:I ANALOG_POL:I
*.PININFO ANALOG_SEL:I ENABLE_VDDA_H:I ENABLE_VSWITCH_H:I HLD_I_H_N:I
*.PININFO NGA_PAD_VPMP_H:O NGB_PAD_VPMP_H:O NGHS_H:I OUT:I PAD:B
*.PININFO PD_CSD_H:O PGHS_H:I PU_CSD_H:O PUG_H[1]:B PUG_H[0]:B VCCD:I
*.PININFO VDDA:I VDDIO:I VDDIO_Q:I VPB_DRVR:B VSSA:I VSSD:I VSSIO:I
*.PININFO VSWITCH:I
XI78 HLD_I_H_N hld_i_h_amux_sw VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
XBBM_logic ANALOG_EN ANALOG_POL ANALOG_SEL ENABLE_VDDA_H enable_vdda_h_n
+ ENABLE_VSWITCH_H HLD_I_H_N nga_amx_vpmp_h NGA_PAD_VPMP_H ngb_amx_vpmp_h
+ NGB_PAD_VPMP_H nmida_vccd nmidb_vccd OUT PD_CSD_H pga_amx_vdda_h_n
+ pga_pad_vddioq_h_n pgb_amx_vdda_h_n pgb_pad_vddioq_h_n PU_CSD_H VCCD VDDA
+ VDDIO_Q VSSA VSSD VSWITCH sky130_fd_io__gpiov2_amux_ctl_logic_i2c_fix
xI77 VSSA VDDA sky130_fd_io__condiode
XI26 net128 net142 sky130_fd_io__res75only_small
XI58 net126 net139 sky130_fd_io__res75only_small
XI28 net124 net144 sky130_fd_io__res75only_small
XI57 PAD net126 sky130_fd_io__res75only_small
XI27 net120 net143 sky130_fd_io__res75only_small
XI55 PAD net128 sky130_fd_io__res75only_small
XI54 PAD net124 sky130_fd_io__res75only_small
XI53 PAD net120 sky130_fd_io__res75only_small
Xmux_a_q0 AMUXBUS_A nga_amx_vpmp_h NGA_PAD_VPMP_H NGHS_H nmida_vccd net144
+ net144 net139 net139 net143 net142 enable_vdda_h_n hld_i_h_amux_sw
+ pga_amx_vdda_h_n pga_pad_vddioq_h_n PGHS_H PUG_H[0] VDDA VDDIO VPB_DRVR VSSA
+ VSSD VSSIO sky130_fd_io__gpio_ovtv2_amux_switch
Xmux_b_q0 AMUXBUS_B ngb_amx_vpmp_h NGB_PAD_VPMP_H NGHS_H nmidb_vccd net144
+ net144 net139 net139 net143 net142 enable_vdda_h_n hld_i_h_amux_sw
+ pgb_amx_vdda_h_n pgb_pad_vddioq_h_n PGHS_H PUG_H[1] VDDA VDDIO VPB_DRVR VSSA
+ VSSD VSSIO sky130_fd_io__gpio_ovtv2_amux_switch
.ENDS sky130_fd_io__gpio_ovtv2_amux_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_amux_switch AG_HV NG_AG_VPMP NG_PAD_VPMP NGHS_H
+ NMID_VDDA PAD_HV_N0 PAD_HV_N1 PAD_HV_N2 PAD_HV_N3 PAD_HV_P0 PAD_HV_P1 PD_H_VDDA
+ PD_H_VDDIO PG_AG_VDDA PG_PAD_VDDIOQ PGHS_H PUG_H VDDA VDDIO VPB_DRVR VSSA VSSD
+ VSSIO
*.PININFO AG_HV:B NG_AG_VPMP:I NG_PAD_VPMP:I NGHS_H:I NMID_VDDA:I
*.PININFO PAD_HV_N0:B PAD_HV_N1:B PAD_HV_N2:B PAD_HV_N3:B PAD_HV_P0:B
*.PININFO PAD_HV_P1:B PD_H_VDDA:I PD_H_VDDIO:I PG_AG_VDDA:I
*.PININFO PG_PAD_VDDIOQ:I PGHS_H:I PUG_H:B VDDA:I VDDIO:I VPB_DRVR:B
*.PININFO VSSA:I VSSD:I VSSIO:I
xI72 VSSA VDDIO sky130_fd_io__condiode
xI71 mid1 VDDIO sky130_fd_io__condiode
xI70 mid VDDIO sky130_fd_io__condiode
XI56 VSSA net85 sky130_fd_io__res75only_small
XI12 VSSA net83 sky130_fd_io__res75only_small
XI46 PAD_HV_N3 NG_PAD_VPMP mid1 mid1 sky130_fd_pr__nfet_g5v0d10v5 m=2 w=10.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI35 mid NG_PAD_VPMP PAD_HV_N1 mid sky130_fd_pr__nfet_g5v0d10v5 m=2 w=10.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI24 PAD_HV_N0 NG_PAD_VPMP mid mid sky130_fd_pr__nfet_g5v0d10v5 m=3 w=10.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI45 mid1 NG_PAD_VPMP PAD_HV_N2 mid1 sky130_fd_pr__nfet_g5v0d10v5 m=3 w=10.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI28 mid NG_AG_VPMP AG_HV mid sky130_fd_pr__nfet_g5v0d10v5 m=5 w=10.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI57 mid1 NMID_VDDA net85 VSSA sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI63 PUG_H NGHS_H PG_PAD_VDDIOQ VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI47 mid1 NG_AG_VPMP AG_HV mid1 sky130_fd_pr__nfet_g5v0d10v5 m=5 w=10.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI75<1> mid PD_H_VDDA VSSA net050<0> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI75<0> mid1 PD_H_VDDA VSSA net050<1> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI74<1> mid PD_H_VDDIO VSSA net051<0> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI74<0> mid1 PD_H_VDDIO VSSA net051<1> sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 mid NMID_VDDA net83 VSSA sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI22 mid PUG_H PAD_HV_P1 VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=10.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI36 mid PUG_H PAD_HV_P0 VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=10.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI62 PG_PAD_VDDIOQ PGHS_H PUG_H VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI26 mid PG_AG_VDDA AG_HV VDDA sky130_fd_pr__pfet_g5v0d10v5 m=4 w=10.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_amux_switch

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

* Modified by Tim to add the additional pin on signal_5_sym_hv_local_5term
* needed to represent the connection from the end of the annular m1 resistor
* (short) back to VDDIO_Q

.SUBCKT sky130_fd_io__gpio_ovtv2_buf_localesd IN_H OUT_H OUT_VT VDDIO_Q VSSD
+ VTRIP_SEL_H
*.PININFO IN_H:I OUT_H:O OUT_VT:O VDDIO_Q:B VSSD:B VTRIP_SEL_H:I
Xesd_res_q0 IN_H OUT_H sky130_fd_io__res250only_small
Xggnfet6_q0 VSSD VDDIO_Q VSSD VDDIO_Q OUT_H VDDIO_Q
+ sky130_fd_io__signal_5_sym_hv_local_5term
Xggnfet1_q0 VSSD OUT_H VSSD VDDIO_Q VSSD VDDIO_Q
+ sky130_fd_io__signal_5_sym_hv_local_5term
Xhv_passgate_q0 OUT_H VTRIP_SEL_H OUT_VT VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=3.0 l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_buf_localesd

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_ctl_hld_i2c_fix ENABLE_H HLD_H_N HLD_I_H_N
+ HLD_I_OVR_H HLD_OVR OD_I_H_N VCC_IO VGND VPWR
*.PININFO ENABLE_H:I HLD_H_N:I HLD_I_H_N:O HLD_I_OVR_H:O HLD_OVR:I
*.PININFO OD_I_H_N:O VCC_IO:I VGND:I VPWR:I
Xhld_nand_q0 ENABLE_H HLD_H_N n1 VGND VCC_IO sky130_fd_io__enh_nand2_1_sp
XI50 OD_I_H_N net45 VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
XI46 n1 n1 n2 VGND VCC_IO sky130_fd_io__enh_nor2_x1
XI49 od_h od_h OD_I_H_N VGND VCC_IO sky130_fd_io__enh_nor2_x1
XI48 ENABLE_H ENABLE_H od_h VGND VCC_IO sky130_fd_io__enh_nand2_1
XI155 n3 n3 HLD_I_H_N VGND VCC_IO sky130_fd_io__nor2_4_enhpath
XI154 n2 n2 n3 VGND VCC_IO sky130_fd_io__nand2_2_enhpath
Xhld_ovr_ls_q0 n2 HLD_OVR hld_ovr_h net79 od_h VGND VCC_IO VGND VPWR
+ sky130_fd_io__com_ctl_ls
XI30 net45 hld_i_ovr_h_n HLD_I_OVR_H VGND VCC_IO sky130_fd_io__hvsbt_nor
XI26 n2 hld_ovr_h hld_i_ovr_h_n VGND VCC_IO sky130_fd_io__hvsbt_nor
.ENDS sky130_fd_io__gpio_ovtv2_ctl_hld_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_ctl_lsbank_i2c_fix DM[2] DM[1] DM[0] DM_H[2]
+ DM_H[1] DM_H[0] DM_H_N[2] DM_H_N[1] DM_H_N[0] HLD_I_H_N HYST_TRIM HYST_TRIM_H
+ HYST_TRIM_H_N IB_MODE_SEL[1] IB_MODE_SEL[0] IB_MODE_SEL_H[1] IB_MODE_SEL_H[0]
+ IB_MODE_SEL_H_N[1] IB_MODE_SEL_H_N[0] INP_DIS INP_DIS_H INP_DIS_H_N OD_I_H_N
+ SLEW_CTL[1] SLEW_CTL[0] SLEW_CTL_H[1] SLEW_CTL_H[0] SLEW_CTL_H_N[1]
+ SLEW_CTL_H_N[0] STARTUP_RST_H STARTUP_ST_H VCC_IO VGND VPWR VTRIP_SEL
+ VTRIP_SEL_H VTRIP_SEL_H_N
*.PININFO DM[2]:I DM[1]:I DM[0]:I DM_H[2]:O DM_H[1]:O DM_H[0]:O
*.PININFO DM_H_N[2]:O DM_H_N[1]:O DM_H_N[0]:O HLD_I_H_N:I HYST_TRIM:I
*.PININFO HYST_TRIM_H:O HYST_TRIM_H_N:O IB_MODE_SEL[1]:I
*.PININFO IB_MODE_SEL[0]:I IB_MODE_SEL_H[1]:O IB_MODE_SEL_H[0]:O
*.PININFO IB_MODE_SEL_H_N[1]:O IB_MODE_SEL_H_N[0]:O INP_DIS:I
*.PININFO INP_DIS_H:O INP_DIS_H_N:O OD_I_H_N:I SLEW_CTL[1]:I
*.PININFO SLEW_CTL[0]:I SLEW_CTL_H[1]:O SLEW_CTL_H[0]:O
*.PININFO SLEW_CTL_H_N[1]:O SLEW_CTL_H_N[0]:O STARTUP_RST_H:I
*.PININFO STARTUP_ST_H:I VCC_IO:I VGND:I VPWR:I VTRIP_SEL:I
*.PININFO VTRIP_SEL_H:O VTRIP_SEL_H_N:O
XI836 OD_I_H_N od_i_h VGND VCC_IO sky130_fd_io__hvsbt_inv_x2
Xtrip_sel_st_q0 trip_sel_st_h od_i_h VGND sky130_fd_io__tk_opti
XI803<1> dm_st_h<1> od_i_h VGND sky130_fd_io__tk_opti
Xtrip_sel_rst_q0 trip_sel_rst_h VGND od_i_h sky130_fd_io__tk_opti
XI802<1> dm_st_h<2> od_i_h VGND sky130_fd_io__tk_opti
XI804<1> dm_rst_h<2> VGND od_i_h sky130_fd_io__tk_opti
XI338<1> dm_rst_h<0> STARTUP_ST_H STARTUP_RST_H sky130_fd_io__tk_opti
XI615 hyst_trim_st_h od_i_h VGND sky130_fd_io__tk_opti
XI614 hyst_trim_rst_h VGND od_i_h sky130_fd_io__tk_opti
XI598<1> ib_mode_sel_st_h<1> od_i_h VGND sky130_fd_io__tk_opti
XI598<0> ib_mode_sel_st_h<0> od_i_h VGND sky130_fd_io__tk_opti
XI597<1> ib_mode_sel_rst_h<1> VGND od_i_h sky130_fd_io__tk_opti
XI597<0> ib_mode_sel_rst_h<0> VGND od_i_h sky130_fd_io__tk_opti
XI337<1> dm_st_h<0> STARTUP_RST_H STARTUP_ST_H sky130_fd_io__tk_opti
XI805<1> dm_rst_h<1> VGND od_i_h sky130_fd_io__tk_opti
XI666<1> slew_ctl_st_h<1> od_i_h VGND sky130_fd_io__tk_opti
XI666<0> slew_ctl_st_h<0> od_i_h VGND sky130_fd_io__tk_opti
XI665<1> slew_ctl_rst_h<1> VGND od_i_h sky130_fd_io__tk_opti
XI665<0> slew_ctl_rst_h<0> VGND od_i_h sky130_fd_io__tk_opti
XI687 ie_n_st_h STARTUP_ST_H STARTUP_RST_H sky130_fd_io__tk_opti
XI686 ie_n_rst_h STARTUP_RST_H STARTUP_ST_H sky130_fd_io__tk_opti
Xdm_ls_0_q0 HLD_I_H_N DM[0] DM_H[0] DM_H_N[0] dm_rst_h<0> dm_st_h<0> VCC_IO VGND
+ VPWR sky130_fd_io__com_ctl_ls
Xinp_dis_ls_q0 HLD_I_H_N INP_DIS INP_DIS_H INP_DIS_H_N ie_n_rst_h ie_n_st_h
+ VCC_IO VGND VPWR sky130_fd_io__com_ctl_ls
Xtrip_sel_ls_q0 HLD_I_H_N VTRIP_SEL VTRIP_SEL_H VTRIP_SEL_H_N trip_sel_rst_h
+ trip_sel_st_h VCC_IO VGND VPWR sky130_fd_io__com_ctl_ls
XI616 HLD_I_H_N HYST_TRIM HYST_TRIM_H HYST_TRIM_H_N hyst_trim_rst_h
+ hyst_trim_st_h VCC_IO VGND VPWR sky130_fd_io__com_ctl_ls
XI595<1> HLD_I_H_N IB_MODE_SEL[1] IB_MODE_SEL_H[1] IB_MODE_SEL_H_N[1]
+ ib_mode_sel_rst_h<1> ib_mode_sel_st_h<1> net58<0> net56<0> net57<0>
+ sky130_fd_io__com_ctl_ls
XI595<0> HLD_I_H_N IB_MODE_SEL[0] IB_MODE_SEL_H[0] IB_MODE_SEL_H_N[0]
+ ib_mode_sel_rst_h<0> ib_mode_sel_st_h<0> net58<1> net56<1> net57<1>
+ sky130_fd_io__com_ctl_ls
XI667<1> HLD_I_H_N SLEW_CTL[1] SLEW_CTL_H[1] SLEW_CTL_H_N[1] slew_ctl_rst_h<1>
+ slew_ctl_st_h<1> net61<0> net59<0> net60<0> sky130_fd_io__com_ctl_ls
XI667<0> HLD_I_H_N SLEW_CTL[0] SLEW_CTL_H[0] SLEW_CTL_H_N[0] slew_ctl_rst_h<0>
+ slew_ctl_st_h<0> net61<1> net59<1> net60<1> sky130_fd_io__com_ctl_ls
Xdm_ls<2>_q0 HLD_I_H_N DM[2] DM_H[2] DM_H_N[2] dm_rst_h<2> dm_st_h<2> VCC_IO
+ VGND VPWR sky130_fd_io__com_ctl_ls
Xdm_ls<1>_q0 HLD_I_H_N DM[1] DM_H[1] DM_H_N[1] dm_rst_h<1> dm_st_h<1> VCC_IO
+ VGND VPWR sky130_fd_io__com_ctl_ls
.ENDS sky130_fd_io__gpio_ovtv2_ctl_lsbank_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_bias PSWG_H VCC_IO VPB_DRVR
*.PININFO PSWG_H:I VCC_IO:I VPB_DRVR:O
Xpsw_vccio_q0 VPB_DRVR PSWG_H VCC_IO VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=22
+ w=15.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI36 VPB_DRVR PSWG_H VCC_IO VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=9 w=10.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_hotswap_bias

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_ctl_i2c_fix EN_H ENHS_LAT_H_N
+ FORCEHI_H[1] OD_I_H_N P3OUT PAD_ESD PGHS_H VDDIO VPB_DRVR VPWR_KA VSSD
*.PININFO EN_H:I ENHS_LAT_H_N:O FORCEHI_H[1]:I OD_I_H_N:I P3OUT:O
*.PININFO PAD_ESD:I PGHS_H:B VDDIO:I VPB_DRVR:I VPWR_KA:I VSSD:I
Xhslog_q0 dishs_h dishs_h_n EN_H enhs_h enhs_h_n enhs_lathys_h_n exiths_h
+ FORCEHI_H[1] OD_I_H_N VDDIO VSSD sky130_fd_io__sio_hotswap_log_i2c_fix
Xhslatch_q0 dishs_h dishs_h_n enhs_h enhs_h_n ENHS_LAT_H_N enhs_lathys_h_n
+ exiths_h P3OUT PAD_ESD PGHS_H VDDIO VSSD VPB_DRVR VPWR_KA
+ sky130_fd_io__gpio_ovtv2_hotswap_latch
.ENDS sky130_fd_io__gpio_ovtv2_hotswap_ctl_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_i2c_fix_leak_fix FORCE_H[1] NGHS_H
+ OD_I_H_N OE_HS_H P2G PAD PAD_ESD PGHS_H PUG_H[7] PUG_H[6] PUG_H[5] PUG_H[4]
+ PUG_H[3] PUG_H[2] PUG_H[1] PUG_H[0] VCC_IO_SOFT VDDIO VPB_DRVR VPWR_KA VSSD
*.PININFO FORCE_H[1]:I NGHS_H:O OD_I_H_N:I OE_HS_H:I P2G:O PAD:I
*.PININFO PAD_ESD:I PGHS_H:O PUG_H[7]:B PUG_H[6]:B PUG_H[5]:B
*.PININFO PUG_H[4]:B PUG_H[3]:B PUG_H[2]:B PUG_H[1]:B PUG_H[0]:B
*.PININFO VCC_IO_SOFT:O VDDIO:I VPB_DRVR:O VPWR_KA:I VSSD:I
Xnon_overlap_q0 p1g NGHS_H P2G padlo VSSD VPB_DRVR
+ sky130_fd_io__gpio_ovtv2_hotswap_nonoverlap_leak_fix
Xpug47_q0 padlo PUG_H[4] PUG_H[7] tie_hi VPB_DRVR
+ sky130_fd_io__gpio_ovtv2_hotswap_pug_ovtfix
Xpghs_q0 OE_HS_H FORCE_H[1] OD_I_H_N net74 PAD_ESD padlo p1g tie_hi VCC_IO_SOFT
+ VDDIO VPB_DRVR VPWR_KA VSSD sky130_fd_io__gpio_ovtv2_hotswap_pghs_i2c_fix
Xresd_tiehi_q0 VPB_DRVR tie_hi sky130_fd_io__sio_tk_tie_r_out_esd
Xresd_vccio_q0 VDDIO VCC_IO_SOFT sky130_fd_io__sio_tk_tie_r_out_esd
Xpug<3>_q0 PAD_ESD padlo PUG_H[3] tie_hi VPB_DRVR
+ sky130_fd_io__gpio_ovtv2_hotswap_pug
Xpug<2>_q0 PAD_ESD padlo PUG_H[2] tie_hi VPB_DRVR
+ sky130_fd_io__gpio_ovtv2_hotswap_pug
Xpug<1>_q0 PAD_ESD padlo PUG_H[1] tie_hi VPB_DRVR
+ sky130_fd_io__gpio_ovtv2_hotswap_pug
Xpug<0>_q0 PAD_ESD padlo PUG_H[0] tie_hi VPB_DRVR
+ sky130_fd_io__gpio_ovtv2_hotswap_pug
Xpug<6>_q0 PAD_ESD padlo PUG_H[6] tie_hi VPB_DRVR
+ sky130_fd_io__gpio_ovtv2_hotswap_pug
Xpug<5>_q0 PAD_ESD padlo PUG_H[5] tie_hi VPB_DRVR
+ sky130_fd_io__gpio_ovtv2_hotswap_pug
Xp1_bias_q0 p1g VDDIO VPB_DRVR sky130_fd_io__gpio_ovtv2_hotswap_bias
Xp2p4_bias_q0 P2G PAD VCC_IO_SOFT VCC_IO_SOFT VPB_DRVR
+ sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias
RI26 P2G net137 short
RI39 P2G net74 short
RI49 PGHS_H p1g short
.ENDS sky130_fd_io__gpio_ovtv2_hotswap_i2c_fix_leak_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_latch DISHS_H DISHS_H_N ENHS_H ENHS_H_N
+ ENHS_LAT_H_N ENHS_LATHYS_H_N EXITHS_H P3OUT PAD_ESD PGHS_H VCC_IO VGND VPB_DRVR
+ VPWR_KA
*.PININFO DISHS_H:I DISHS_H_N:I ENHS_H:I ENHS_H_N:I ENHS_LAT_H_N:O
*.PININFO ENHS_LATHYS_H_N:O EXITHS_H:I P3OUT:O PAD_ESD:I PGHS_H:B
*.PININFO VCC_IO:I VGND:I VPB_DRVR:I VPWR_KA:I
XI660 VGND net102 VGND VGND VCC_IO VCC_IO sky130_fd_io__sio_hvsbt_inv_x1
XI528 n6 net96 VGND VGND VCC_IO VCC_IO sky130_fd_io__sio_hvsbt_inv_x1
XEhys2 ENHS_LATHYS_H_N ENHS_LAT_H_N sky130_fd_io__tk_em1o
XI658 net96 ENHS_LAT_H_N sky130_fd_io__tk_em1s
XEhys1 net117 ENHS_LATHYS_H_N sky130_fd_io__tk_em1s
Xhys_q0 n6 net117 VCC_IO VGND sky130_fd_io__sio_hotswap_hys
Xpghspd_q0 ENHS_H n2 PGHS_H VGND sky130_fd_io__sio_hotswap_pghspd
Xwpdenhs_q0 VPWR_KA net127 VGND sky130_fd_io__sio_hotswap_wpd
Xwpdexhs_q0 VPWR_KA net124 VGND sky130_fd_io__sio_hotswap_wpd
XI502 net186 PGHS_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI484 net161 ENHS_H PGHS_H VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI491 n5 n6 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI498 n2 n6 net124 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI500 net170 ENHS_H_N n2 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xnexiths_q0 PGHS_H EXITHS_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI485 n3 n2 net161 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI499 n4 PGHS_H net170 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI497 n6 n5 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xndishs_q0 PGHS_H DISHS_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI508 n2 ENHS_H_N net186 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI696 VGND EXITHS_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI487 PGHS_H n5 net127 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI697 VGND DISHS_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI492 n5 n6 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI503 n4 VGND VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=2.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI488 n3 VGND VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=2.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI505 n6 n5 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI493 n5 n3 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI323 n2 DISHS_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=4 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI279 n2 PAD_ESD VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=4 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI504 n6 n4 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI689 P3OUT PAD_ESD VCC_IO VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=12 w=10.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_hotswap_latch

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_nonoverlap_leak_fix P1G P1GB P2G PADLO
+ VGND VPWR
*.PININFO P1G:O P1GB:O P2G:O PADLO:I VGND:I VPWR:I
XI76 P1G P1GB VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI64 p1g_new PADLO VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI53 padlo_bar PADLO VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI50 p2g_new p1g_new VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI49 p2g_new padlo_bar VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI65 p1g_new p2g_new VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI77 P2G p2gb VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI70 p2gb p2g_new VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI72 P1GB p1g_new VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI54 padlo_bar PADLO VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI69 p1g_new PADLO net140 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=4.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI78 P2G p2gb VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=0.42 l=2.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI67 net140 p2g_new VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=8.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI71 p2gb p2g_new VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI79 P1G P1GB VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=2.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI51 p2g_new padlo_bar net124 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=4.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI73 P1GB p1g_new VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI52 net124 p1g_new VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=8.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_hotswap_nonoverlap_leak_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_pghs_i2c_fix EN_H FORCE_H[1] OD_I_H_N
+ P3OUT PAD PADLO PGHS_H TIE_HI VCC_IO_SOFT VDDIO VPB_DRVR VPWR_KA VSSD
*.PININFO EN_H:I FORCE_H[1]:I OD_I_H_N:I P3OUT:O PAD:I PADLO:O
*.PININFO PGHS_H:O TIE_HI:I VCC_IO_SOFT:I VDDIO:I VPB_DRVR:I VPWR_KA:I
*.PININFO VSSD:I
Xhsctl_q0 EN_H enhs_lat_h_n FORCE_H[1] OD_I_H_N P3OUT PAD net50 VDDIO VPB_DRVR
+ VPWR_KA VSSD sky130_fd_io__gpio_ovtv2_hotswap_ctl_i2c_fix
XI3 enhs_latbuf_h_n PADLO sky130_fd_io__sio_tk_em1s
XEpghs12 PGHS_H net54 sky130_fd_io__sio_tk_em1o
XI2 enhs_lat_h enhs_latbuf_h_n VSSD VSSD VDDIO VDDIO
+ sky130_fd_io__sio_hvsbt_inv_x4
XI1 enhs_lat_h_n enhs_lat_h VSSD VSSD VDDIO VDDIO sky130_fd_io__sio_hvsbt_inv_x1
Xpghspu_q0 PAD PGHS_H net50 TIE_HI VCC_IO_SOFT VPB_DRVR
+ sky130_fd_io__gpio_ovtv2_hotswap_pghspu
Xclamp_q0 VSSD VDDIO VSSD VDDIO PAD VDDIO sky130_fd_io__signal_5_sym_hv_local_5term
Xpghs12_q0 net54 PADLO VPB_DRVR VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0
+ l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_hotswap_pghs_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_pghspu PAD PGHS_H PGHS_H_LATCH TIE_HI
+ VCC_IO_SOFT VPB_DRVR
*.PININFO PAD:I PGHS_H:O PGHS_H_LATCH:O TIE_HI:I VCC_IO_SOFT:I
*.PININFO VPB_DRVR:I
XEg9 TIE_HI pg8 sky130_fd_io__sio_tk_em1o
XEg2 pg2 VCC_IO_SOFT sky130_fd_io__sio_tk_em1s
XEg5 pg6 pg4 sky130_fd_io__sio_tk_em1s
XEg4 pg4 pg3 sky130_fd_io__sio_tk_em1s
XEpghs3 padhi3 PGHS_H_LATCH sky130_fd_io__sio_tk_em1s
XEg3 pg3 pg2 sky130_fd_io__sio_tk_em1s
XEpghs7 padhi7 net36 sky130_fd_io__sio_tk_em1s
XEg7 pg7 pg6 sky130_fd_io__sio_tk_em1s
XEg8 pg8 pg7 sky130_fd_io__sio_tk_em1s
XEpghs2 padhi2 padhi3 sky130_fd_io__sio_tk_em1s
XEpghs8 PGHS_H padhi7 sky130_fd_io__sio_tk_em1s
Xpghs8_q0 PGHS_H pg8 PAD VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=20.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xpghs2_q0 padhi2 pg2 PAD VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=20.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xpghs3_q0 padhi3 pg3 PAD VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=20.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xpghs6_q0 net36 pg6 PAD VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=15.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xpghs4_q0 PGHS_H_LATCH pg4 PAD VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=15.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xpghs7_q0 padhi7 pg7 PAD VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=20.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_hotswap_pghspu

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_pug PAD PADLO PUG_H TIE_HI VPB_DRVR
*.PININFO PAD:I PADLO:I PUG_H:O TIE_HI:I VPB_DRVR:I
XEg1 PADLO net22 sky130_fd_io__sio_tk_em1s
XI65 net24 TIE_HI sky130_fd_io__sio_tk_em1s
XEs2 net26 TIE_HI sky130_fd_io__sio_tk_em1s
XEs1 PAD net26 sky130_fd_io__sio_tk_em1o
XEg2 net22 net24 sky130_fd_io__sio_tk_em1o
XI52 PUG_H net22 net26 VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=15.0 l=0.5
+ mult=1 sa=1.825 sb=1.825 sd=0.28 topography=normal area=0.063 perim=1.14
XI53 PUG_H net24 net26 VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=15.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_hotswap_pug

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_pug_ovtfix PADLO PUG4_H PUG7_H TIE_HI
+ VPB_DRVR
*.PININFO PADLO:I PUG4_H:O PUG7_H:O TIE_HI:I VPB_DRVR:I
XI52 PUG4_H PADLO TIE_HI VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=15.0 l=0.5
+ mult=1 sa=1.825 sb=1.825 sd=0.28 topography=normal area=0.063 perim=1.14
XI53 PUG7_H PADLO TIE_HI VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=15.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_hotswap_pug_ovtfix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias P2G PAD SOFT_VCC_IO TIE_HI
+ VPB_DRVR
*.PININFO P2G:I PAD:I SOFT_VCC_IO:I TIE_HI:I VPB_DRVR:B
Xpsw_pad4_q0 VPB_DRVR VPB_DRVR P2G PAD
+ sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit
Xpsw_pad0_q0 VPB_DRVR VPB_DRVR P2G PAD
+ sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit
Xpsw_pad3_q0 VPB_DRVR VPB_DRVR P2G PAD
+ sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit
Xpsw_pad2_q0 VPB_DRVR VPB_DRVR P2G PAD
+ sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit
Xpsw_pad5_q0 VPB_DRVR VPB_DRVR SOFT_VCC_IO PAD
+ sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit
Xpsw_pad1_q0 VPB_DRVR VPB_DRVR P2G PAD
+ sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit
XI5 TIE_HI SOFT_VCC_IO sky130_fd_io__tk_em1o
.ENDS sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit PB PD PGIN PS
*.PININFO PB:I PD:B PGIN:I PS:B
Xpdrv_q0 PD PGIN PS PB sky130_fd_pr__esd_pfet_g5v0d10v5 m=2 w=15.5 l=0.55 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_ibuf_se EN_H EN_H_N ENABLE_VDDIO_LV IBUFMUX_OUT
+ IBUFMUX_OUT_H IN_H IN_VT MODE_NORMAL_N MODE_REF_3V_N MODE_REF_N MODE_VCCD_N
+ VCCHIB VDDIO_Q VREFIN VSSD VTRIP_SEL_H VTRIP_SEL_H_N
*.PININFO EN_H:I EN_H_N:I ENABLE_VDDIO_LV:I IBUFMUX_OUT:O
*.PININFO IBUFMUX_OUT_H:O IN_H:I IN_VT:I MODE_NORMAL_N:I
*.PININFO MODE_REF_3V_N:I MODE_REF_N:I MODE_VCCD_N:I VCCHIB:I
*.PININFO VDDIO_Q:I VREFIN:I VSSD:I VTRIP_SEL_H:I VTRIP_SEL_H_N:I
Xlvls_q0 ENABLE_VDDIO_LV out IBUFMUX_OUT net43 VCCHIB VSSD
+ sky130_fd_io__gpio_ovtv2_ipath_lvls
Xhvls_q0 EN_H_N out out_n IBUFMUX_OUT_H net49 VDDIO_Q VSSD
+ sky130_fd_io__gpio_ovtv2_ipath_hvls
Xbuf_q0 EN_H EN_H_N ENABLE_VDDIO_LV IN_H IN_VT MODE_NORMAL_N MODE_REF_3V_N
+ MODE_REF_N MODE_VCCD_N out out_n VCCHIB VDDIO_Q VREFIN VSSD VTRIP_SEL_H
+ VTRIP_SEL_H_N sky130_fd_io__gpio_ovtv2_in_buf
.ENDS sky130_fd_io__gpio_ovtv2_ibuf_se

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_ictl_logic DM_H_N[2] DM_H_N[1] DM_H_N[0]
+ HYS_TRIM IBUF_MODE_SEL[0] IBUF_MODE_SEL[1] INP_DIS_H_N INP_DIS_I_H INP_DIS_I_H_N
+ MODE_NORMAL_N MODE_REF_3V_N MODE_REF_N MODE_VCCD_N TRIPSEL_I_H TRIPSEL_I_H_N
+ VDDIO_Q VSSD VTRIP_SEL_H
*.PININFO DM_H_N[2]:I DM_H_N[1]:I DM_H_N[0]:I HYS_TRIM:I
*.PININFO IBUF_MODE_SEL[0]:I IBUF_MODE_SEL[1]:I INP_DIS_H_N:I
*.PININFO INP_DIS_I_H:O INP_DIS_I_H_N:O MODE_NORMAL_N:O
*.PININFO MODE_REF_3V_N:O MODE_REF_N:O MODE_VCCD_N:O TRIPSEL_I_H:O
*.PININFO TRIPSEL_I_H_N:O VDDIO_Q:I VSSD:I VTRIP_SEL_H:I
XI41 net66 MODE_NORMAL_N TRIPSEL_I_H VSSD VDDIO_Q sky130_fd_io__hvsbt_nor
XI34 IBUF_MODE_SEL[1] net70 net60 VSSD VDDIO_Q sky130_fd_io__hvsbt_nor
XI33 IBUF_MODE_SEL[1] IBUF_MODE_SEL[0] net55 VSSD VDDIO_Q
+ sky130_fd_io__hvsbt_nor
Xdm10nand_inv_q0 nand_dm01 and_dm01 VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
XI68 INP_DIS_I_H INP_DIS_I_H_N VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
XI43 TRIPSEL_I_H TRIPSEL_I_H_N VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
XI50 MODE_REF_N mode_ref VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
XI39 IBUF_MODE_SEL[0] net70 VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
XI61 VTRIP_SEL_H net66 VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
Xinpdis_q0 dm_buf_dis INP_DIS_H_N INP_DIS_I_H VSSD VDDIO_Q
+ sky130_fd_io__hvsbt_nand2
Xdm210_q0 DM_H_N[2] and_dm01 dm_buf_dis VSSD VDDIO_Q sky130_fd_io__hvsbt_nand2
Xdm10_q0 DM_H_N[1] DM_H_N[0] nand_dm01 VSSD VDDIO_Q sky130_fd_io__hvsbt_nand2
XI40 INP_DIS_I_H_N IBUF_MODE_SEL[1] MODE_REF_N VSSD VDDIO_Q
+ sky130_fd_io__hvsbt_nand2
XI36 INP_DIS_I_H_N net60 MODE_VCCD_N VSSD VDDIO_Q sky130_fd_io__hvsbt_nand2
XI35 INP_DIS_I_H_N net55 MODE_NORMAL_N VSSD VDDIO_Q sky130_fd_io__hvsbt_nand2
XI52 mode_ref HYS_TRIM MODE_REF_3V_N VSSD VDDIO_Q sky130_fd_io__hvsbt_nand2
.ENDS sky130_fd_io__gpio_ovtv2_ictl_logic

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_in_buf EN_H EN_H_N ENABLE_VDDIO_LV IN_H IN_VT
+ MODE_NORMAL_N MODE_REF_3V_N MODE_REF_N MODE_VCCD_N OUT OUT_N VCCHIB VDDIO_Q
+ VREFIN VSSD VTRIP_SEL_H VTRIP_SEL_H_N
*.PININFO EN_H:I EN_H_N:I ENABLE_VDDIO_LV:I IN_H:I IN_VT:I
*.PININFO MODE_NORMAL_N:I MODE_REF_3V_N:I MODE_REF_N:I MODE_VCCD_N:I
*.PININFO OUT:O OUT_N:O VCCHIB:I VDDIO_Q:I VREFIN:I VSSD:I
*.PININFO VTRIP_SEL_H:I VTRIP_SEL_H_N:I
XI35 ENABLE_VDDIO_LV EN_H enable_vddio_lv_n VSSD VCCHIB
+ sky130_fd_io__hvsbt_nand2
xI405 virt_pwr1 VDDIO_Q sky130_fd_io__condiode
xI404 virt_pwr VDDIO_Q sky130_fd_io__condiode
XI488 VTRIP_SEL_H MODE_NORMAL_N mode_normal_cmos_h VSSD VDDIO_Q
+ sky130_fd_io__hvsbt_nor
XI43 mode_normal_cmos_h mode_normal_cmos_h_n VSSD VDDIO_Q
+ sky130_fd_io__hvsbt_inv_x1
XI630 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI105 fbk1 in_b fbk VSSD sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI620 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI441 IN_VT VTRIP_SEL_H_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI417 OUT EN_H_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI419 OUT_N EN_H_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI394 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI494 fbk IN_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=6 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 fbk2 in_b fbk VSSD sky130_fd_pr__nfet_g5v0d10v5 m=3 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI26 OUT in_b VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI49 vddio_ref VREFIN virt_pwr virt_pwr sky130_fd_pr__nfet_05v0_nvt m=3 w=10.0
+ l=0.9 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI451 fbk IN_VT VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=12 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI453 in_b IN_H fbk VSSD sky130_fd_pr__nfet_g5v0d10v5 m=6 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI111 vddio_ref1 VREFIN virt_pwr1 virt_pwr1 sky130_fd_pr__nfet_05v0_nvt m=3
+ w=10.0 l=0.9 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI446 OUT_N OUT VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI389 virt_pwr VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0 l=0.8
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI450 in_b IN_VT fbk VSSD sky130_fd_pr__nfet_g5v0d10v5 m=6 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI274 fbk1 MODE_REF_N virt_pwr1 virt_pwr1 sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI116 virt_pwr MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=2
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI109 in_b IN_H virt_pwr virt_pwr sky130_fd_pr__pfet_g5v0d10v5 m=3 w=5.0 l=0.8
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI25 OUT in_b virt_pwr1 virt_pwr1 sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI13 fbk2 mode_normal_cmos_h_n VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=2
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI611 fbk1 MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI396 vddio_ref1 MODE_REF_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=2
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI115 virt_pwr MODE_VCCD_N vcchib_int virt_pwr sky130_fd_pr__pfet_g5v0d10v5 m=4
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI478 vcchib_int1 enable_vddio_lv_n VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 m=8
+ w=5.0 l=0.25 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI373 vddio_ref MODE_REF_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=2
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI403 OUT in_b virt_pwr2 virt_pwr2 sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI376 fbk2 MODE_REF_3V_N virt_pwr1 virt_pwr1 sky130_fd_pr__pfet_g5v0d10v5 m=4
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI477 vcchib_int enable_vddio_lv_n VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 m=8
+ w=5.0 l=0.25 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI401 in_b IN_H virt_pwr2 virt_pwr2 sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.8
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI457 OUT_N OUT virt_pwr1 virt_pwr1 sky130_fd_pr__pfet_g5v0d10v5 m=5 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI486 fbk1 MODE_VCCD_N vcchib_int virt_pwr1 sky130_fd_pr__pfet_g5v0d10v5 m=2
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI400 virt_pwr2 MODE_VCCD_N vcchib_int virt_pwr2 sky130_fd_pr__pfet_g5v0d10v5
+ m=2 w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI381 virt_pwr1 MODE_VCCD_N vcchib_int1 virt_pwr1 sky130_fd_pr__pfet_g5v0d10v5
+ m=6 w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI380 virt_pwr1 MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=2
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_in_buf

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_ipath DM_H_N[2] DM_H_N[1] DM_H_N[0]
+ ENABLE_VDDIO_LV HYS_TRIM_H IB_MODE_SEL_H[1] IB_MODE_SEL_H[0] INP_DIS_H_N OUT
+ OUT_H PAD VCCHIB VDDIO_Q VINREF VSSD VTRIP_SEL_H
*.PININFO DM_H_N[2]:I DM_H_N[1]:I DM_H_N[0]:I ENABLE_VDDIO_LV:I
*.PININFO HYS_TRIM_H:I IB_MODE_SEL_H[1]:I IB_MODE_SEL_H[0]:I
*.PININFO INP_DIS_H_N:I OUT:O OUT_H:O PAD:B VCCHIB:I VDDIO_Q:I
*.PININFO VINREF:B VSSD:I VTRIP_SEL_H:I
Xibuf_se_q0 en_h en_h_n ENABLE_VDDIO_LV OUT OUT_H in_h in_vt mode_normal_n
+ mode_ref_3v_n mode_ref_n mode_vccd_n VCCHIB VDDIO_Q VINREF VSSD tripsel_i_h
+ tripsel_i_h_n sky130_fd_io__gpio_ovtv2_ibuf_se
Xesd_q0 PAD in_h in_vt VDDIO_Q VSSD tripsel_i_h
+ sky130_fd_io__gpio_ovtv2_buf_localesd
Xlogic_q0 DM_H_N[2] DM_H_N[1] DM_H_N[0] HYS_TRIM_H IB_MODE_SEL_H[0]
+ IB_MODE_SEL_H[1] INP_DIS_H_N en_h_n en_h mode_normal_n mode_ref_3v_n mode_ref_n
+ mode_vccd_n tripsel_i_h tripsel_i_h_n VDDIO_Q VSSD VTRIP_SEL_H
+ sky130_fd_io__gpio_ovtv2_ictl_logic
.ENDS sky130_fd_io__gpio_ovtv2_ipath

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_ipath_hvls EN_H_N IN INB OUT OUT_B VDDIO_Q VSSD
*.PININFO EN_H_N:I IN:I INB:I OUT:O OUT_B:O VDDIO_Q:I VSSD:I
XI250 fbk fbk_b VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI253 OUT OUT_B VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=5 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI249 fbk_b fbk VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI248 OUT_B fbk VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI247 OUT_B fbk VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI252 OUT OUT_B VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=3 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI304 fbk INB VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=3 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI262 fbk EN_H_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI246 fbk_b IN VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=3 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_ipath_hvls

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_ipath_lvls ENABLE_VDDIO_LV IN OUT OUT_B VCCHIB
+ VSSD
*.PININFO ENABLE_VDDIO_LV:I IN:I OUT:O OUT_B:O VCCHIB:I VSSD:I
XI248 fbk_n IN VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI271 OUT OUT_B VCCHIB VCCHIB sky130_fd_pr__pfet_01v8_hvt m=2 w=5.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI281 fbk_n ENABLE_VDDIO_LV VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI272 OUT_B fbk VCCHIB VCCHIB sky130_fd_pr__pfet_01v8_hvt m=1 w=5.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI277 fbk fbk_n VCCHIB VCCHIB sky130_fd_pr__pfet_01v8_hvt m=1 w=5.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI273 OUT OUT_B VSSD VSSD sky130_fd_pr__nfet_01v8 m=2 w=3.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI278 fbk fbk_n VSSD VSSD sky130_fd_pr__nfet_01v8 m=1 w=3.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI305 OUT_B fbk VSSD VSSD sky130_fd_pr__nfet_01v8 m=1 w=3.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI535 fbk_n IN vssd_1 VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI279 vssd_1 ENABLE_VDDIO_LV VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_ipath_lvls

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_obpredrvr_leak_fix DRVHI_H DRVLO_H_N
+ I2C_MODE_H_N NGHS_H OE_I_H_N PAD PD_DIS_H PD_H[3] PD_H[2] PD_H[1] PD_H[0]
+ PDEN_H_N[1] PDEN_H_N[0] PGHS_H PU_H_N[3] PU_H_N[2] PU_H_N[1] PU_H_N[0] PUEN_H[1]
+ PUEN_H[0] PUG_H SLEW_CTL_H[1] SLEW_CTL_H[0] SLEW_CTL_H_N[1] SLEW_CTL_H_N[0]
+ SLOW_H SLOW_H_N VCC_IO VGND_IO VPB_DRVR VSSD
*.PININFO DRVHI_H:I DRVLO_H_N:I I2C_MODE_H_N:I NGHS_H:I OE_I_H_N:I
*.PININFO PAD:B PD_DIS_H:I PD_H[3]:O PD_H[2]:O PD_H[1]:O PD_H[0]:O
*.PININFO PDEN_H_N[1]:I PDEN_H_N[0]:I PGHS_H:I PU_H_N[3]:O PU_H_N[2]:O
*.PININFO PU_H_N[1]:O PU_H_N[0]:O PUEN_H[1]:I PUEN_H[0]:I PUG_H:I
*.PININFO SLEW_CTL_H[1]:I SLEW_CTL_H[0]:I SLEW_CTL_H_N[1]:I
*.PININFO SLEW_CTL_H_N[0]:I SLOW_H:I SLOW_H_N:I VCC_IO:I VGND_IO:I
*.PININFO VPB_DRVR:I VSSD:I
XI192 DRVLO_H_N en_cmos_b I2C_MODE_H_N NGHS_H nsw_en OE_I_H_N PAD PD_DIS_H
+ PD_H[3] PD_H[2] PDEN_H_N[1] PGHS_H PUG_H SLEW_CTL_H[1] SLEW_CTL_H[0]
+ SLEW_CTL_H_N[1] SLEW_CTL_H_N[0] SLOW_H_N VCC_IO VGND_IO VPB_DRVR VSSD
+ sky130_fd_io__gpio_ovtv2_obpredrvr_new_leak_fix
XI191 DRVHI_H DRVLO_H_N en_cmos_b nsw_en PD_H[3] PD_H[2] PD_H[1] PD_H[0]
+ PDEN_H_N[1] PDEN_H_N[0] PU_H_N[3] PU_H_N[2] PU_H_N[1] PU_H_N[0] PUEN_H[1]
+ PUEN_H[0] SLOW_H SLOW_H_N VCC_IO VGND_IO sky130_fd_io__gpio_ovtv2_obpredrvr_old
.ENDS sky130_fd_io__gpio_ovtv2_obpredrvr_leak_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_obpredrvr_new_leak_fix DRVLO_H_N EN_CMOS_B
+ I2C_MODE_H_N NGHS_H NSW_EN OE_I_H_N PAD PD_DIS_H PD_H[3] PD_H[2] PDEN_H_N[1]
+ PGHS_H PUG_H SLEW_CTL_H[1] SLEW_CTL_H[0] SLEW_CTL_H_N[1] SLEW_CTL_H_N[0]
+ SLOW_H_N VCC_IO VGND_IO VPB_DRVR VSSD
*.PININFO DRVLO_H_N:I EN_CMOS_B:O I2C_MODE_H_N:I NGHS_H:I NSW_EN:O
*.PININFO OE_I_H_N:I PAD:B PD_DIS_H:I PD_H[3]:O PD_H[2]:O
*.PININFO PDEN_H_N[1]:I PGHS_H:I PUG_H:I SLEW_CTL_H[1]:I
*.PININFO SLEW_CTL_H[0]:I SLEW_CTL_H_N[1]:I SLEW_CTL_H_N[0]:I
*.PININFO SLOW_H_N:I VCC_IO:I VGND_IO:I VPB_DRVR:I VSSD:I
Xpd_strong_q0 DRVLO_H_N EN_CMOS_B I2C_MODE_H_N NGHS_H NSW_EN OE_I_H_N PAD
+ PD_DIS_H PD_H[3] PD_H[2] PDEN_H_N[1] PGHS_H PUG_H SLEW_CTL_H[1] SLEW_CTL_H[0]
+ SLEW_CTL_H_N[1] SLEW_CTL_H_N[0] SLOW_H_N VCC_IO VGND_IO VPB_DRVR VSSD
+ sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_leak_fix
.ENDS sky130_fd_io__gpio_ovtv2_obpredrvr_new_leak_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_obpredrvr_old DRVHI_H DRVLO_H_N EN_CMOS_B
+ NSW_EN PD_H[3] PD_H[2] PD_H[1] PD_H[0] PDEN_H_N[1] PDEN_H_N[0] PU_H_N[3]
+ PU_H_N[2] PU_H_N[1] PU_H_N[0] PUEN_H[1] PUEN_H[0] SLOW_H SLOW_H_N VCC_IO VGND_IO
*.PININFO DRVHI_H:I DRVLO_H_N:I EN_CMOS_B:I NSW_EN:I PD_H[3]:O
*.PININFO PD_H[2]:O PD_H[1]:O PD_H[0]:O PDEN_H_N[1]:I PDEN_H_N[0]:I
*.PININFO PU_H_N[3]:O PU_H_N[2]:O PU_H_N[1]:O PU_H_N[0]:O PUEN_H[1]:I
*.PININFO PUEN_H[0]:I SLOW_H:I SLOW_H_N:I VCC_IO:I VGND_IO:I
xI19 VGND_IO VCC_IO sky130_fd_io__condiode
Xpu_strong_slow_q0 DRVHI_H PU_H_N[1] PUEN_H[1] VCC_IO VGND_IO
+ sky130_fd_io__com_pupredrvr_strong_slow
Xpu_weak_q0 DRVHI_H PU_H_N[0] PUEN_H[0] VCC_IO VGND_IO
+ sky130_fd_io__com_pupredrvr_weak
XI151 DRVLO_H_N PD_H[0] PDEN_H_N[0] VCC_IO VGND_IO
+ sky130_fd_io__com_pdpredrvr_weak
Xpd_strong_slow_q0 DRVLO_H_N PD_H[1] EN_CMOS_B VCC_IO VGND_IO
+ sky130_fd_io__com_pdpredrvr_strong_slow
XI150 DRVLO_H_N DRVLO_H_N EN_CMOS_B NSW_EN PD_H[3] PD_H[2] PDEN_H_N[1] SLOW_H
+ VCC_IO VGND_IO sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_cmos
Xpu_strong_q0 DRVHI_H PU_H_N[3] PU_H_N[2] PUEN_H[1] SLOW_H_N VCC_IO VGND_IO
+ sky130_fd_io__gpio_ovtv2_pupredrvr_strong
.ENDS sky130_fd_io__gpio_ovtv2_obpredrvr_old

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_octl_dat_i2c_fix_leak_fix DM_H[2] DM_H[1]
+ DM_H[0] DM_H_N[2] DM_H_N[1] DM_H_N[0] DRVHI_H HLD_I_H_N HLD_I_OVR_H NGHS_H
+ OD_I_H_N OE_HS_H OE_N OUT PAD PD_H[3] PD_H[2] PD_H[1] PD_H[0] PGHS_H PU_H_N[3]
+ PU_H_N[2] PU_H_N[1] PU_H_N[0] PUG_H SLEW_CTL_H[1] SLEW_CTL_H[0] SLEW_CTL_H_N[1]
+ SLEW_CTL_H_N[0] SLOW SLOW_H_N VCCD VDDIO VPB_DRVR VPWR_KA VSSD VSSIO
*.PININFO DM_H[2]:I DM_H[1]:I DM_H[0]:I DM_H_N[2]:I DM_H_N[1]:I
*.PININFO DM_H_N[0]:I DRVHI_H:O HLD_I_H_N:I HLD_I_OVR_H:I NGHS_H:I
*.PININFO OD_I_H_N:I OE_HS_H:O OE_N:I OUT:I PAD:B PD_H[3]:O PD_H[2]:O
*.PININFO PD_H[1]:O PD_H[0]:O PGHS_H:I PU_H_N[3]:O PU_H_N[2]:O
*.PININFO PU_H_N[1]:O PU_H_N[0]:O PUG_H:I SLEW_CTL_H[1]:I
*.PININFO SLEW_CTL_H[0]:I SLEW_CTL_H_N[1]:I SLEW_CTL_H_N[0]:I SLOW:I
*.PININFO SLOW_H_N:O VCCD:I VDDIO:I VPB_DRVR:I VPWR_KA:I VSSD:I
*.PININFO VSSIO:I
Xpredrvr_q0 DRVHI_H drvlo_h_n pden_h_n<2> NGHS_H oe_i_h_n PAD net72 PD_H[3]
+ PD_H[2] PD_H[1] PD_H[0] pden_h_n<1> pden_h_n<0> PGHS_H PU_H_N[3] PU_H_N[2]
+ PU_H_N[1] PU_H_N[0] puen_h<1> puen_h<0> PUG_H SLEW_CTL_H[1] SLEW_CTL_H[0]
+ SLEW_CTL_H_N[1] SLEW_CTL_H_N[0] slow_h SLOW_H_N VDDIO VSSIO VPB_DRVR VSSD
+ sky130_fd_io__gpio_ovtv2_obpredrvr_leak_fix
Xdatoe_q0 DRVHI_H drvlo_h_n HLD_I_H_N HLD_I_OVR_H OD_I_H_N oe_h OE_N OUT net72
+ VDDIO VSSD VPWR_KA sky130_fd_io__gpio_ovtv2_opath_datoe_i2c_fix
Xctl_q0 DM_H[2] DM_H[1] DM_H[0] DM_H_N[2] DM_H_N[1] DM_H_N[0] HLD_I_H_N OD_I_H_N
+ pden_h_n<2> pden_h_n<1> pden_h_n<0> net86 net85 puen_h<1> puen_h<0> SLOW slow_h
+ SLOW_H_N VDDIO VSSD VCCD VDDIO sky130_fd_io__gpio_ovtv2_octl_i2c_fix
XI354 oe_hs_i_h oe_hs_i_h_n VSSD VSSD VDDIO VDDIO sky130_fd_io__sio_hvsbt_inv_x1
XI353 oe_h oe_i_h_n VSSD VSSD VDDIO VDDIO sky130_fd_io__sio_hvsbt_inv_x2
XI355 oe_hs_i_h_n OE_HS_H VSSD VSSD VDDIO VDDIO sky130_fd_io__sio_hvsbt_inv_x2
XI351 net86 net85 n<1> VSSD VSSD VDDIO VDDIO sky130_fd_io__sio_hvsbt_nor
XI352 n<1> oe_i_h_n oe_hs_i_h VSSD VSSD VDDIO VDDIO sky130_fd_io__sio_hvsbt_nor
.ENDS sky130_fd_io__gpio_ovtv2_octl_dat_i2c_fix_leak_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_octl_i2c_fix DM_H[2] DM_H[1] DM_H[0] DM_H_N[2]
+ DM_H_N[1] DM_H_N[0] HLD_I_H_N OD_I_H_N PDEN_H_N[2] PDEN_H_N[1] PDEN_H_N[0]
+ PUEN_0_H PUEN_2OR1_H PUEN_H[1] PUEN_H[0] SLOW SLOW_H SLOW_H_N VCC_IO VGND VPWR
+ VREG_EN_H_N
*.PININFO DM_H[2]:I DM_H[1]:I DM_H[0]:I DM_H_N[2]:I DM_H_N[1]:I
*.PININFO DM_H_N[0]:I HLD_I_H_N:I OD_I_H_N:I PDEN_H_N[2]:O
*.PININFO PDEN_H_N[1]:O PDEN_H_N[0]:O PUEN_0_H:O PUEN_2OR1_H:O
*.PININFO PUEN_H[1]:O PUEN_H[0]:O SLOW:I SLOW_H:O SLOW_H_N:O VCC_IO:I
*.PININFO VGND:I VPWR:I VREG_EN_H_N:I
XI211 n<8> DM_H_N[1] PUEN_0_H VGND VCC_IO sky130_fd_io__hvsbt_nor
XI201 DM_H_N[2] DM_H_N[1] n<9> VGND VCC_IO sky130_fd_io__hvsbt_nor
XI366 DM_H[1] DM_H[0] net87 VGND VCC_IO sky130_fd_io__hvsbt_nor
XI210 DM_H[2] DM_H[0] n<8> VGND VCC_IO sky130_fd_io__hvsbt_xor
XI200 DM_H[2] DM_H[1] n<10> VGND VCC_IO sky130_fd_io__hvsbt_xor
XI185 DM_H_N[0] n<4> net207 VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI186 DM_H_N[2] DM_H_N[1] n<4> VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI187 DM_H[1] DM_H[0] n<3> VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI208 PUEN_2OR1_H VREG_EN_H_N n<5> VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI203 n<10> DM_H[0] n<1> VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI204 n<9> DM_H_N[0] n<0> VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI205 n<1> n<0> PUEN_2OR1_H VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI365 net87 DM_H[2] PDEN_H_N[2] VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI254 puen_h1_n PUEN_H[1] VGND VCC_IO sky130_fd_io__hvsbt_inv_x2
XI256 puen_h0_n PUEN_H[0] VGND VCC_IO sky130_fd_io__hvsbt_inv_x2
XI249 pden_h0 PDEN_H_N[0] VGND VCC_IO sky130_fd_io__hvsbt_inv_x2
XI247 pden_h1 PDEN_H_N[1] VGND VCC_IO sky130_fd_io__hvsbt_inv_x2
XI377 PUEN_0_H puen_h0_n VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
XI209 n<5> n<2> VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
XI376 n<2> puen_h1_n VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
XI374 net207 pden_h1 VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
XI375 n<3> pden_h0 VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
XI381 OD_I_H_N n9 VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
Xls_slow_q0 HLD_I_H_N SLOW SLOW_H SLOW_H_N n9 VGND VCC_IO VGND VPWR
+ sky130_fd_io__com_ctl_ls
.ENDS sky130_fd_io__gpio_ovtv2_octl_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_odrvr_i2c_fix_leak_fix FORCE_H[1]
+ NGA_PAD_VPMP_H NGB_PAD_VPMP_H NGHS_H OD_I_H_N OE_HS_H PAD PD_CSD_H PD_H[3]
+ PD_H[2] PD_H[1] PD_H[0] PGHS_H PU_CSD_H PU_H_N[3] PU_H_N[2] PU_H_N[1] PU_H_N[0]
+ PUG_H[7] PUG_H[6] PUG_H[5] TIE_HI_ESD TIE_LO_ESD VDDIO VDDIO_AMX VPB_DRVR VSSA
+ VSSD VSSIO VSSIO_AMX
*.PININFO FORCE_H[1]:I NGA_PAD_VPMP_H:I NGB_PAD_VPMP_H:I NGHS_H:O
*.PININFO OD_I_H_N:I OE_HS_H:I PAD:O PD_CSD_H:I PD_H[3]:I PD_H[2]:I
*.PININFO PD_H[1]:I PD_H[0]:I PGHS_H:O PU_CSD_H:I PU_H_N[3]:I
*.PININFO PU_H_N[2]:I PU_H_N[1]:I PU_H_N[0]:I PUG_H[7]:B PUG_H[6]:B
*.PININFO PUG_H[5]:B TIE_HI_ESD:O TIE_LO_ESD:O VDDIO:I VDDIO_AMX:B
*.PININFO VPB_DRVR:B VSSA:I VSSD:I VSSIO:I VSSIO_AMX:I
Xhotswap_q0 FORCE_H[1] NGHS_H OD_I_H_N OE_HS_H p2g PAD pad_esd PGHS_H PUG_H[7]
+ PUG_H[6] PUG_H[5] pug_h<4> pug_h<3> pug_h<2> pug_h<1> pug_h<0> net74 VDDIO
+ VPB_DRVR VDDIO VSSD sky130_fd_io__gpio_ovtv2_hotswap_i2c_fix_leak_fix
Xbondpad_q0 PAD VSSIO sky130_fd_io__com_pad
Xodrvr_q0 TIE_HI_ESD PAD pad_esd PD_CSD_H PD_H[3] PD_H[2] PD_H[1] PD_H[0] PGHS_H
+ PU_CSD_H PU_H_N[3] PU_H_N[2] PU_H_N[1] PU_H_N[0] pug_h<4> pug_h<3> pug_h<2>
+ pug_h<1> pug_h<0> TIE_HI_ESD TIE_LO_ESD VDDIO VDDIO_AMX VPB_DRVR VSSD VSSIO
+ VSSIO_AMX sky130_fd_io__gpio_ovtv2_odrvr_sub
XI122<2> PD_H[3] PGHS_H net106<0> VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI122<1> PD_H[2] PGHS_H net106<1> VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI122<0> PD_H[1] PGHS_H net106<2> VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI85<2> net106<0> PGHS_H VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI85<1> net106<1> PGHS_H VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI85<0> net106<2> PGHS_H VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI104<2> net102<0> PGHS_H VSSA VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI104<1> net102<1> PGHS_H VSSA VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI104<0> net102<2> PGHS_H VSSA VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI103<2> PD_CSD_H PGHS_H net102<0> VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI103<1> NGA_PAD_VPMP_H PGHS_H net102<1> VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=0.42 l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI103<0> NGB_PAD_VPMP_H PGHS_H net102<2> VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=0.42 l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_odrvr_i2c_fix_leak_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_odrvr_sub NGHS_H PAD PAD_ESD PD_CSD_H PD_H[3]
+ PD_H[2] PD_H[1] PD_H[0] PGHS_H PU_CSD_H PU_H_N[3] PU_H_N[2] PU_H_N[1] PU_H_N[0]
+ PUG_H[4] PUG_H[3] PUG_H[2] PUG_H[1] PUG_H[0] TIE_HI_ESD TIE_LO_ESD VDDIO
+ VDDIO_AMX VPB_DRVR VSSD VSSIO VSSIO_AMX
*.PININFO NGHS_H:I PAD:B PAD_ESD:B PD_CSD_H:I PD_H[3]:I PD_H[2]:I
*.PININFO PD_H[1]:I PD_H[0]:I PGHS_H:I PU_CSD_H:I PU_H_N[3]:I
*.PININFO PU_H_N[2]:I PU_H_N[1]:I PU_H_N[0]:I PUG_H[4]:B PUG_H[3]:B
*.PININFO PUG_H[2]:B PUG_H[1]:B PUG_H[0]:B TIE_HI_ESD:B TIE_LO_ESD:B
*.PININFO VDDIO:I VDDIO_AMX:B VPB_DRVR:B VSSD:I VSSIO:I VSSIO_AMX:I
Xpddrvr_strong_slow_q0 strong_slow_pad PD_H[1] VDDIO VSSIO
+ sky130_fd_io__gpio_pddrvr_strong_slow
XI73 weak_pad PD_H[0] VDDIO VSSIO sky130_fd_io__gpio_pddrvr_weak
Xres_q0 strong_slow_pad PAD_ESD VSSIO sky130_fd_io__com_res_strong_slow
Xres_weak_q0 weak_pad PAD_ESD VSSIO sky130_fd_io__com_res_weak
Xpd_drvr_q0 PAD PD_CSD_H PD_H[3] PD_H[2] TIE_LO_ESD VDDIO VSSIO VSSIO_AMX
+ sky130_fd_io__gpio_ovtv2_pddrvr
Xpudrvr_weak_q0 NGHS_H weak_pad PGHS_H PU_H_N[0] PUG_H[0] VDDIO VPB_DRVR VSSD
+ VSSIO sky130_fd_io__gpio_ovtv2_pudrvr_weak
Xstrong_slow_pudrvr_q0 NGHS_H strong_slow_pad PGHS_H PU_H_N[1] PUG_H[1] VDDIO
+ VPB_DRVR VSSD VSSIO sky130_fd_io__gpio_ovtv2_pudrvr_strong_slow
Xpudrvr_strong_q0 NGHS_H NGHS_H NGHS_H PAD PGHS_H PGHS_H PGHS_H PU_CSD_H
+ PU_H_N[3] PU_H_N[2] PUG_H[4] PUG_H[3] PUG_H[2] TIE_HI_ESD VDDIO VDDIO_AMX
+ VPB_DRVR VSSD VSSIO sky130_fd_io__gpio_ovtv2_pudrvr_strong
Xres_esd_q0 PAD_ESD PAD sky130_fd_io__res75only_small
xI72 VSSIO VDDIO sky130_fd_io__condiode
.ENDS sky130_fd_io__gpio_ovtv2_odrvr_sub

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_opath_datoe_i2c_fix DRVHI_H DRVLO_H_N HLD_H_N
+ HLD_I_OVR_H OD_I_H_N OE_H OE_N OUT PD_DIS_H VCC_IO VGND VPWR_KA
*.PININFO DRVHI_H:O DRVLO_H_N:O HLD_H_N:I HLD_I_OVR_H:I OD_I_H_N:I
*.PININFO OE_H:O OE_N:I OUT:I PD_DIS_H:O VCC_IO:I VGND:I VPWR_KA:I
Xdat_ls_q0 HLD_I_OVR_H OUT PD_DIS_H pu_dis_h VGND net60 VCC_IO VGND VPWR_KA
+ sky130_fd_io__gpio_dat_ls
Xcclat_q0 DRVHI_H DRVLO_H_N OE_H PD_DIS_H pu_dis_h VCC_IO VGND
+ sky130_fd_io__com_cclat_i2c_fix
XI36 OD_I_H_N net60 VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
XI37 OD_I_H_N net56 VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
Xoe_ls_q0 HLD_I_OVR_H OE_N OE_H net56 OD_I_H_N VCC_IO VGND VPWR_KA
+ sky130_fd_io__gpio_dat_ls_i2c_fix
.ENDS sky130_fd_io__gpio_ovtv2_opath_datoe_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_opath_i2c_fix_leak_fix DM_H[2] DM_H[1] DM_H[0]
+ DM_H_N[2] DM_H_N[1] DM_H_N[0] HLD_I_H_N HLD_I_OVR_H NGA_PAD_VPMP_H
+ NGB_PAD_VPMP_H OD_I_H_N OE_N OUT PAD PD_CSD_H PGHS_H PU_CSD_H PUG_H[6] PUG_H[5]
+ SLEW_CTL_H[1] SLEW_CTL_H[0] SLEW_CTL_H_N[1] SLEW_CTL_H_N[0] SLOW TIE_HI_ESD
+ TIE_LO_ESD VCCD VDDIO VDDIO_AMX VPB_DRVR VPWR_KA VSSA VSSD VSSIO VSSIO_AMX
*.PININFO DM_H[2]:I DM_H[1]:I DM_H[0]:I DM_H_N[2]:I DM_H_N[1]:I
*.PININFO DM_H_N[0]:I HLD_I_H_N:I HLD_I_OVR_H:I NGA_PAD_VPMP_H:I
*.PININFO NGB_PAD_VPMP_H:I OD_I_H_N:I OE_N:I OUT:I PAD:O PD_CSD_H:I
*.PININFO PGHS_H:O PU_CSD_H:I PUG_H[6]:B PUG_H[5]:B SLEW_CTL_H[1]:I
*.PININFO SLEW_CTL_H[0]:I SLEW_CTL_H_N[1]:I SLEW_CTL_H_N[0]:I SLOW:I
*.PININFO TIE_HI_ESD:O TIE_LO_ESD:O VCCD:I VDDIO:I VDDIO_AMX:B
*.PININFO VPB_DRVR:B VPWR_KA:I VSSA:I VSSD:I VSSIO:I VSSIO_AMX:I
Xodrvr_q0 TIE_LO_ESD NGA_PAD_VPMP_H NGB_PAD_VPMP_H nghs_h OD_I_H_N oe_hs_h PAD
+ PD_CSD_H pd_h<3> pd_h<2> pd_h<1> pd_h<0> PGHS_H PU_CSD_H pu_h_n<3> pu_h_n<2>
+ pu_h_n<1> pu_h_n<0> pug_h<7> PUG_H[6] PUG_H[5] TIE_HI_ESD TIE_LO_ESD VDDIO
+ VDDIO_AMX VPB_DRVR VSSA VSSD VSSIO VSSIO_AMX
+ sky130_fd_io__gpio_ovtv2_odrvr_i2c_fix_leak_fix
Xopath_q0 DM_H[2] DM_H[1] DM_H[0] DM_H_N[2] DM_H_N[1] DM_H_N[0] drvhi_h
+ HLD_I_H_N HLD_I_OVR_H nghs_h OD_I_H_N oe_hs_h OE_N OUT PAD pd_h<3> pd_h<2>
+ pd_h<1> pd_h<0> PGHS_H pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> pug_h<7>
+ SLEW_CTL_H[1] SLEW_CTL_H[0] SLEW_CTL_H_N[1] SLEW_CTL_H_N[0] SLOW slow_h_n VCCD
+ VDDIO VPB_DRVR VPWR_KA VSSD VSSIO
+ sky130_fd_io__gpio_ovtv2_octl_dat_i2c_fix_leak_fix
.ENDS sky130_fd_io__gpio_ovtv2_opath_i2c_fix_leak_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_pddrvr PAD PD_CSD PD_H[3] PD_H[2] TIE_LO_ESD
+ VDDIO VSSIO VSSIO_Q
*.PININFO PAD:B PD_CSD:I PD_H[3]:I PD_H[2]:I TIE_LO_ESD:O VDDIO:B
*.PININFO VSSIO:B VSSIO_Q:B
XI26 VSSIO TIE_LO_ESD sky130_fd_io__tk_tie_r_out_esd
Xn1_q0 PAD PD_H[2] VSSIO sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn2_q0 PAD PD_H[2] VSSIO sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn3_q0 PAD PD_H[2] VSSIO sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn8_q0 PAD PD_H[3] VSSIO sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn7_q0 PAD PD_H[3] VSSIO sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn6_q0 PAD PD_H[3] VSSIO sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn5_q0 PAD PD_H[3] VSSIO sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn9_q0 PAD PD_H[3] VSSIO sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn10_q0 PAD PD_H[3] VSSIO sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn11_q0 PAD PD_H[3] VSSIO sky130_fd_io__gpio_ovtv2_pddrvr_unit
xI9 VSSIO VDDIO sky130_fd_io__condiode
xI62 VSSIO_Q VDDIO sky130_fd_io__condiode
RI8 VDDIO net96 short
Xn14_q0 PAD PD_CSD VSSIO_Q VSSIO_Q sky130_fd_pr__esd_nfet_g5v0d10v5 m=1 w=40.31
+ l=0.55 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xn13_q0 PAD PD_CSD VSSIO_Q VSSIO_Q sky130_fd_pr__esd_nfet_g5v0d10v5 m=1 w=40.31
+ l=0.55 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_pddrvr

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_pddrvr_unit ND NGIN NS
*.PININFO ND:B NGIN:I NS:B
Xndrv_q0 ND NGIN NS NS sky130_fd_pr__esd_nfet_g5v0d10v5 m=1 w=40.31 l=0.55
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_pddrvr_unit

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_pdpredrvr_pbias DRVLO_H_N EN_H EN_H_N PBIAS
+ PD_H PDEN_H_N VCC_IO VGND_IO
*.PININFO DRVLO_H_N:I EN_H:I EN_H_N:I PBIAS:O PD_H:I PDEN_H_N:I
*.PININFO VCC_IO:I VGND_IO:I
XE1 n<1> n<0> sky130_fd_io__tk_em1o
XE2 PBIAS pbias1 sky130_fd_io__tk_em1o
XE3 pbias1 net88 sky130_fd_io__tk_em1s
XE4 net108 PBIAS sky130_fd_io__tk_em1s
XE6 PBIAS net84 sky130_fd_io__tk_em1s
XE5 n<101> bias_g sky130_fd_io__tk_em1s
XI27 n<0> PD_H EN_H_N sky130_fd_io__tk_opto
XI47 PBIAS bias_g VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.0 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI24 n<1> DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI18 bias_g DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI23 n<0> n<0> n<1> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI13 drvlo_i_h DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI20 bias_g n<1> VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI19 bias_g EN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI34 net157 bias_g VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI36 net108 bias_g VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.0 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI38 n<1> PDEN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI48 n<100> PD_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=4.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI41 n<101> PD_H n<100> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=4.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI44 PBIAS PBIAS pbias1 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=8 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI45 pbias1 pbias1 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=8 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI15 net183 EN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=10.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI16 net171 n<0> net183 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=10.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 PBIAS EN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 drvlo_i_h DRVLO_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI17 bias_g DRVLO_H_N net171 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=3 w=7.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI14 PBIAS drvlo_i_h VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI33 N0 VGND_IO VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=8.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI32 net161 net161 N0 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI31 net157 net157 net161 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI30 net88 N0 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=8 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI43 net84 bias_g VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=4.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI40 N0 drvlo_i_h VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_pdpredrvr_pbias

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_cmos DRVHI_H DRVLO_H_N
+ EN_CMOS_B NSW_EN_INT PD_H[3] PD_H[2] PDEN_H_N SLOW_H VCC_IO VGND_IO
*.PININFO DRVHI_H:I DRVLO_H_N:I EN_CMOS_B:I NSW_EN_INT:I PD_H[3]:O
*.PININFO PD_H[2]:O PDEN_H_N:I SLOW_H:I VCC_IO:I VGND_IO:I
Xbias_q0 DRVHI_H en_fast_h en_fast_h_n pbias_out PD_H[2] PDEN_H_N VCC_IO VGND_IO
+ sky130_fd_io__gpio_ovtv2_pdpredrvr_pbias
Xnr3_q0 DRVLO_H_N net76 net76 PD_H[2] NSW_EN_INT VCC_IO VGND_IO
+ sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_nr2
Xnr2_q0 DRVLO_H_N en_fast2_n<1> en_fast2_n<0> PD_H[3] NSW_EN_INT VCC_IO VGND_IO
+ sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_nr3
XI77 en_fast2_n<1> pbias_out en_fast_h_n sky130_fd_io__tk_opto
XI76 net76 pbias_out en_fast_h_n sky130_fd_io__tk_opto
XI79 en_fast2_n<0> en_fast2_n<1> VCC_IO sky130_fd_io__tk_opti
Xinv_q0 en_fast_h en_fast_h_n VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
Xnor_q0 SLOW_H EN_CMOS_B en_fast_h VGND_IO VCC_IO sky130_fd_io__com_nor2_dnw
.ENDS sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_cmos

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

* Modified by Tim:  Added 3rd terminal to res_generic_nd__hv devices

.SUBCKT sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_leak_fix DRVLO_H_N EN_CMOS_B
+ I2C_MODE_H_N NGHS_H NSW_EN_INT OE_I_H_N PAD_CAP PD_DIS_H PD_H[3] PD_H[2]
+ PDEN_H_N[1] PGHS_H PUG_H SLEW_CTL_H[1] SLEW_CTL_H[0] SLEW_CTL_H_N[1]
+ SLEW_CTL_H_N[0] SLOW_H_N VCC_IO VGND_IO VPB_DRVR VSSD
*.PININFO DRVLO_H_N:I EN_CMOS_B:O I2C_MODE_H_N:I NGHS_H:I NSW_EN_INT:O
*.PININFO OE_I_H_N:I PAD_CAP:B PD_DIS_H:I PD_H[3]:O PD_H[2]:O
*.PININFO PDEN_H_N[1]:I PGHS_H:I PUG_H:I SLEW_CTL_H[1]:I
*.PININFO SLEW_CTL_H[0]:I SLEW_CTL_H_N[1]:I SLEW_CTL_H_N[0]:I
*.PININFO SLOW_H_N:I VCC_IO:I VGND_IO:I VPB_DRVR:I VSSD:I
XI123 PD_DIS_H nsw_enb OE_I_H_N net200 VGND_IO VCC_IO sky130_fd_io__nor3_dnw
xI208 VGND_IO VCC_IO sky130_fd_io__condiode
XI161 net293 drvlo_h_n_i2c_2 VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
XI159 net298 drvlo_h_n_i2c_1 VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
XI224 net288 net247 VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
XI605 en enb VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
XI176 net318 drvlo_h_n_i2c_4 VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
XI191 nsw_en nsw_enb VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
XI198 net303 drvlo_h_n_i2c VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
XI179 net283 NSW_EN_INT VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
XI168 net263 mode1b VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
XI122 drvlo_h drvlo_h_n_buf VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
XI170 net278 mode3b VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
XI715 PDEN_H_N[1] pden_h<1> VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
XI162 net313 drvlo_h_n_i2c_3 VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
XI254 DRVLO_H_N drvlo_h VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
XI602 vdelay net200 en VGND_IO VCC_IO sky130_fd_io__com_nand2_dnw
XI112 pden_h<1> nsw_enb EN_CMOS_B VGND_IO VCC_IO sky130_fd_io__com_nand2_dnw
XI430 SLEW_CTL_H[1] SLEW_CTL_H_N[0] net263 VGND_IO VCC_IO
+ sky130_fd_io__com_nand2_dnw
XI175 drvlo_h_n_i2c mode4b net318 VGND_IO VCC_IO sky130_fd_io__com_nor2_dnw
XI163 drvlo_h_n_i2c mode3b net313 VGND_IO VCC_IO sky130_fd_io__com_nor2_dnw
XI109 SLOW_H_N I2C_MODE_H_N nsw_en VGND_IO VCC_IO sky130_fd_io__com_nor2_dnw
XI197 nsw_enb drvlo_h_n_buf net303 VGND_IO VCC_IO sky130_fd_io__com_nor2_dnw
XI158 drvlo_h_n_i2c mode1b net298 VGND_IO VCC_IO sky130_fd_io__com_nor2_dnw
XI160 drvlo_h_n_i2c mode2b net293 VGND_IO VCC_IO sky130_fd_io__com_nor2_dnw
XI225 SLEW_CTL_H[1] SLEW_CTL_H[0] net288 VGND_IO VCC_IO
+ sky130_fd_io__com_nor2_dnw
XI181 PDEN_H_N[1] nsw_en net283 VGND_IO VCC_IO sky130_fd_io__com_nor2_dnw
XI169 SLEW_CTL_H[1] SLEW_CTL_H_N[0] net278 VGND_IO VCC_IO
+ sky130_fd_io__com_nor2_dnw
XI94 nsw_en nsw_enb PD_H[2] PD_H[3] VCC_IO VGND_IO
+ sky130_fd_io__gpio_ovtv2_predrvr_switch
XI288 N0 net193 VGND_IO sky130_fd_pr__res_generic_nd__hv W=0.5 L=113.375 m=1
XI287 vdiode net190 VGND_IO sky130_fd_pr__res_generic_nd__hv W=0.5 L=113.375 m=1
XI206 N0 en VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI190 net531 en VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI220 net420 enb VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI153 PD_H[2] PDEN_H_N[1] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI182 VGND_IO vdelay VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.0
+ l=2.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI201 net352 N0 net190 VGND_IO sky130_fd_pr__nfet_05v0_nvt m=10 w=1.0 l=0.9
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI625 net404 PD_H[3] net348 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI339 net400 pden_h<1> VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI125 PD_H[3] drvlo_h_n_buf net400 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=4
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI344 PD_H[3] PDEN_H_N[1] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI63 net388 vdiode PD_H[3] VGND_IO sky130_fd_pr__nfet_05v0_nvt m=2 w=10.0 l=0.9
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI189 net388 VGND_IO VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI10 biasp vdiode net336 VGND_IO sky130_fd_pr__nfet_05v0_nvt m=5 w=10.0 l=0.9
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI374 net519 nsw_en PD_H[3] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI137 biasp1 vdiode VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI13 net369 net369 VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=5 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI8 vdiode vdiode VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=5 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI165 vdiode en VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI14 N0 N0 net369 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=5 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI15 net352 N0 net190 VGND_IO sky130_fd_pr__nfet_05v0_nvt m=4 w=10.0 l=0.9
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI755 net348 PD_H[3] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI579 vdelay drvlo_h net404 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI192 net519 VGND_IO VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI219 net336 vdiode vr VGND_IO sky130_fd_pr__nfet_01v8_lvt m=5 w=7.0 l=0.15
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI232<1> cas3 PGHS_H PD_H[3] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI232<0> cas10 PGHS_H PD_H[3] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI278 VGND_IO VGND_IO VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI20 PUG_H NGHS_H nsw_enb VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI245 cas10 VCC_IO cas4 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI196 nc biasp VCC_IO VCC_IO sky130_fd_pr__pfet_01v8 m=5 w=0.55 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI200 cas3 biasp1 nc VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI199 PD_H[3] drvlo_h_n_i2c_2 cas3 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI205 net352 en VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI156 cas5 biasp1 ne VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI580 vdelay drvlo_h VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI136 biasp biasp1 na VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI144 cas4 biasp1 nd VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI84 PD_H[3] drvlo_h_n_i2c cas2 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI230 nc VCC_IO VCC_IO VCC_IO sky130_fd_pr__pfet_01v8 m=1 w=0.55 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI79 nb biasp VCC_IO VCC_IO sky130_fd_pr__pfet_01v8 m=17 w=0.55 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI260 net535 enb VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI228 PD_H[3] drvlo_h_n_i2c net535 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI73 net388 drvlo_h_n_i2c net531 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI561 PD_H[3] drvlo_h_n_i2c_1 cas4 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI560 nd biasp VCC_IO VCC_IO sky130_fd_pr__pfet_01v8 m=14 w=0.55 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI375 PD_H[3] PUG_H net519 VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI164 biasp enb VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI167 biasp1 enb VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI138 biasp1 biasp1 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI145 cas2 biasp1 nb VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI141 na biasp VCC_IO VCC_IO sky130_fd_pr__pfet_01v8 m=10 w=0.55 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI154 ne biasp VCC_IO VCC_IO sky130_fd_pr__pfet_01v8 m=14 w=0.55 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI178 net193 en VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI155 PD_H[3] drvlo_h_n_i2c_3 cas5 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI241 cas10 biasp1 nf VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI240 nf biasp VCC_IO VCC_IO sky130_fd_pr__pfet_01v8 m=8 w=0.55 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI229 ne VCC_IO VCC_IO VCC_IO sky130_fd_pr__pfet_01v8 m=2 w=0.55 l=4.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI217 nb VCC_IO VCC_IO VCC_IO sky130_fd_pr__pfet_01v8 m=3 w=0.55 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI216 nd VCC_IO VCC_IO VCC_IO sky130_fd_pr__pfet_01v8 m=2 w=0.55 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI215 cas3 VCC_IO cas2 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI214 cas5 VCC_IO cas2 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI239 PD_H[3] drvlo_h_n_i2c_3 cas10 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI213 cas3 VCC_IO cas4 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI212 na VCC_IO VCC_IO VCC_IO sky130_fd_pr__pfet_01v8 m=2 w=0.55 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI211 VCC_IO VCC_IO VCC_IO VCC_IO sky130_fd_pr__pfet_01v8 m=4 w=0.55 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI210 VCC_IO VCC_IO VCC_IO VCC_IO sky130_fd_pr__pfet_01v8 m=6 w=0.55 l=4.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI248<5> na enb VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI248<4> nb enb VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI248<3> nc enb VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI248<2> nd enb VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI248<1> ne enb VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI248<0> nf enb VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI30 nsw_enb PGHS_H PUG_H VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI70 net531 en VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
RI221 net420 vr sky130_fd_pr__res_generic_po W=0.75 L=513.445 m=1
RI186 SLEW_CTL_H_N[0] mode4b sky130_fd_pr__res_generic_m1 L=0.035 W=1
RI157 net247 mode2b sky130_fd_pr__res_generic_m1 L=0.035 W=1
.ENDS sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_leak_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_nr2 DRVLO_H_N EN_FAST_N[1]
+ EN_FAST_N[0] PD_H PDEN_H_N VCC_IO VGND_IO
*.PININFO DRVLO_H_N:I EN_FAST_N[1]:I EN_FAST_N[0]:I PD_H:O PDEN_H_N:I
*.PININFO VCC_IO:I VGND_IO:I
Xmnin_q0 PD_H DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=5 w=3.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI56 int_slow PDEN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42
+ l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmpin_slow_q0 PD_H DRVLO_H_N int_slow VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=1.0 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpen_slow_q0 int_slow PDEN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=1.0 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpin_fast<1>_q0 PD_H DRVLO_H_N int_nor<1> net19<0> sky130_fd_pr__pfet_g5v0d10v5
+ m=2 w=3.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpin_fast<0>_q0 PD_H DRVLO_H_N int_nor<0> net19<1> sky130_fd_pr__pfet_g5v0d10v5
+ m=2 w=3.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpen_fast<1>_q0 int_nor<1> EN_FAST_N[1] VCC_IO VCC_IO
+ sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.0 l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xmpen_fast<0>_q0 int_nor<0> EN_FAST_N[0] VCC_IO VCC_IO
+ sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_nr2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_nr3 DRVLO_H_N EN_FAST_N[1]
+ EN_FAST_N[0] PD_H PDEN_H_N VCC_IO VGND_IO
*.PININFO DRVLO_H_N:I EN_FAST_N[1]:I EN_FAST_N[0]:I PD_H:O PDEN_H_N:I
*.PININFO VCC_IO:I VGND_IO:I
Xmnin_q0 PD_H DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=5 w=3.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI56 int_slow PDEN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42
+ l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmpin_slow_q0 PD_H DRVLO_H_N int_slow VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=1.0 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpen_slow_q0 int_slow PDEN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=1.0 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpin_fast<1>_q0 PD_H DRVLO_H_N int_nor<1> net19<0> sky130_fd_pr__pfet_g5v0d10v5
+ m=2 w=3.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpin_fast<0>_q0 PD_H DRVLO_H_N int_nor<0> net19<1> sky130_fd_pr__pfet_g5v0d10v5
+ m=2 w=3.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpen_fast<1>_q0 int_nor<1> EN_FAST_N[1] VCC_IO VCC_IO
+ sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.0 l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xmpen_fast<0>_q0 int_nor<0> EN_FAST_N[0] VCC_IO VCC_IO
+ sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_nr3

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_predrvr_switch NMOS_EN PMOS_EN SIG1 SIG2 VCC_IO
+ VGND_IO
*.PININFO NMOS_EN:I PMOS_EN:I SIG1:B SIG2:B VCC_IO:I VGND_IO:I
XI374 SIG1 NMOS_EN SIG2 VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI375 SIG2 PMOS_EN SIG1 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_predrvr_switch

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_pudrvr_strong NGHS_H[4] NGHS_H[3] NGHS_H[2] PAD
+ PGHS_H[4] PGHS_H[3] PGHS_H[2] PU_CSD_H PU_H_N[3] PU_H_N[2] PUG_H[4] PUG_H[3]
+ PUG_H[2] TIE_HI_ESD VDDIO VDDIO_AMX VPB_DRVR VSSD VSSIO
*.PININFO NGHS_H[4]:I NGHS_H[3]:I NGHS_H[2]:I PAD:B PGHS_H[4]:I
*.PININFO PGHS_H[3]:I PGHS_H[2]:I PU_CSD_H:I PU_H_N[3]:I PU_H_N[2]:I
*.PININFO PUG_H[4]:B PUG_H[3]:B PUG_H[2]:B TIE_HI_ESD:O VDDIO:I
*.PININFO VDDIO_AMX:B VPB_DRVR:B VSSD:I VSSIO:I
XI49 VDDIO TIE_HI_ESD sky130_fd_io__tk_tie_r_out_esd
XI133 VPB_DRVR tie_hi_vpbdrvr sky130_fd_io__tk_tie_r_out_esd
XI112 PUG_H[2] net83 sky130_fd_io__tk_em2o
XI111 PUG_H[4] net81 sky130_fd_io__tk_em2o
XI141 PUG_H[3] net79 sky130_fd_io__tk_em2o
XI152 PUG_H[4] net079 sky130_fd_io__tk_em2o
XI142 tie_hi_vpbdrvr net79 sky130_fd_io__tk_em2s
XI82 tie_hi_vpbdrvr net83 sky130_fd_io__tk_em2s
XI109 tie_hi_vpbdrvr net81 sky130_fd_io__tk_em2s
XI153 tie_hi_vpbdrvr net079 sky130_fd_io__tk_em2s
Xn7_q0 VPB_DRVR PAD PUG_H[3] VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn6_q0 VPB_DRVR PAD PUG_H[3] VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn5<2>_q0 VPB_DRVR PAD PUG_H[3] VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn5<1>_q0 VPB_DRVR PAD PUG_H[3] VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn5<0>_q0 VPB_DRVR PAD PUG_H[3] VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn4_q0 VPB_DRVR PAD PUG_H[2] VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn2<3>_q0 VPB_DRVR PAD net83 VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn2<2>_q0 VPB_DRVR PAD net83 VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn2<1>_q0 VPB_DRVR PAD net83 VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn2<0>_q0 VPB_DRVR PAD net83 VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn9<1>_q0 VPB_DRVR PAD net79 VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn9<0>_q0 VPB_DRVR PAD net79 VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn11<1>_q0 VPB_DRVR PAD PUG_H[4] VDDIO_AMX
+ sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn11<0>_q0 VPB_DRVR PAD PUG_H[4] VDDIO_AMX
+ sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn12<1>_q0 VPB_DRVR PAD net81 VDDIO_AMX sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn12<0>_q0 VPB_DRVR PAD net81 VDDIO_AMX sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn1<1>_q0 VPB_DRVR PAD PUG_H[2] VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn1<0>_q0 VPB_DRVR PAD PUG_H[2] VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn3<1>_q0 VPB_DRVR PAD PUG_H[2] VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn3<0>_q0 VPB_DRVR PAD PUG_H[2] VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn8<1>_q0 VPB_DRVR PAD PUG_H[3] VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn8<0>_q0 VPB_DRVR PAD PUG_H[3] VDDIO sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn10<1>_q0 VPB_DRVR PAD net079 VDDIO_AMX
+ sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn10<0>_q0 VPB_DRVR PAD net079 VDDIO_AMX
+ sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
XI136 PUG_H[4] NGHS_H[4] PU_CSD_H VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI127 PUG_H[2] NGHS_H[2] PU_H_N[2] VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI25 PUG_H[3] NGHS_H[3] PU_H_N[3] VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI137 PU_CSD_H PGHS_H[4] PUG_H[4] VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=2
+ w=3.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI128 PU_H_N[2] PGHS_H[2] PUG_H[2] VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=2
+ w=3.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI24 PU_H_N[3] PGHS_H[3] PUG_H[3] VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=2
+ w=3.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_pudrvr_strong

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_pudrvr_strong_slow NGHS_H PAD PGHS_H PU_H_N
+ PUG_H VDDIO VPB_DRVR VSSD VSSIO
*.PININFO NGHS_H:I PAD:B PGHS_H:I PU_H_N:I PUG_H:B VDDIO:I VPB_DRVR:I
*.PININFO VSSD:I VSSIO:I
XI20 PUG_H NGHS_H PU_H_N VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI30 PU_H_N PGHS_H PUG_H VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xpdrv_q0 PAD PUG_H VDDIO VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=12 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_pudrvr_strong_slow

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5 PB PD PGIN PS
*.PININFO PB:B PD:B PGIN:I PS:B
Xpdrv_q0 PD PGIN PS PB sky130_fd_pr__esd_pfet_g5v0d10v5 m=1 w=15.5 l=0.55 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_pudrvr_weak NGHS_H PAD PGHS_H PU_H_N PUG_H
+ VDDIO VPB_DRVR VSSD VSSIO
*.PININFO NGHS_H:I PAD:B PGHS_H:I PU_H_N:I PUG_H:B VDDIO:I VPB_DRVR:I
*.PININFO VSSD:I VSSIO:I
XI36 PAD net26 sky130_fd_io__tk_em1o
XI51 PUG_H NGHS_H PU_H_N VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI50 PU_H_N PGHS_H PUG_H VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xpdrv_q0 PAD PUG_H VDDIO VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=3 w=10.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI35 net26 PUG_H VDDIO VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=10.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI29 PAD PUG_H VDDIO VPB_DRVR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=10.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_pudrvr_weak

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_pupredrvr_strong DRVHI_H PU_H_N[3] PU_H_N[2]
+ PUEN_H SLOW_H_N VCC_IO VGND_IO
*.PININFO DRVHI_H:I PU_H_N[3]:O PU_H_N[2]:O PUEN_H:I SLOW_H_N:I
*.PININFO VCC_IO:I VGND_IO:I
Xnd2b_q0 DRVHI_H en_fast_h_3<3> en_fast_h_3<2> en_fast_h_3<1> en_fast_h_3<0>
+ PU_H_N[3] PUEN_H VCC_IO VGND_IO sky130_fd_io__gpio_ovtv2_pupredrvr_strong_nd3
Xnd2a_q0 DRVHI_H net54 net54 net54 net54 PU_H_N[2] PUEN_H VCC_IO VGND_IO
+ sky130_fd_io__gpio_ovtv2_pupredrvr_strong_nd2
XI98 en_fast_h_3<0> en_fast_h_3<3> VGND_IO sky130_fd_io__tk_opti
XI97 en_fast_h_3<1> en_fast_h_3<3> VGND_IO sky130_fd_io__tk_opti
XI92 en_fast_h_3<3> nbias_out en_fast_h sky130_fd_io__tk_opto
XI96 en_fast_h_3<2> en_fast_h_3<3> VGND_IO sky130_fd_io__tk_opto
XI93 net54 nbias_out en_fast_h sky130_fd_io__tk_opto
Xinv_q0 en_fast_h_n en_fast_h VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
Xnbias_q0 DRVHI_H en_fast_h en_fast_h_n nbias_out PU_H_N[2] PUEN_H VCC_IO
+ VGND_IO sky130_fd_io__com_pupredrvr_nbias
Xnand_q0 PUEN_H SLOW_H_N en_fast_h_n VGND_IO VCC_IO sky130_fd_io__com_nand2_dnw
.ENDS sky130_fd_io__gpio_ovtv2_pupredrvr_strong

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_pupredrvr_strong_nd2 DRVHI_H EN_FAST[3]
+ EN_FAST[2] EN_FAST[1] EN_FAST[0] PU_H_N PUEN_H VCC_IO VGND_IO
*.PININFO DRVHI_H:I EN_FAST[3]:I EN_FAST[2]:I EN_FAST[1]:I
*.PININFO EN_FAST[0]:I PU_H_N:O PUEN_H:I VCC_IO:I VGND_IO:I
XE1 net30 PU_H_N sky130_fd_io__tk_em1s
Rrespu1 int_res net30 sky130_fd_pr__res_generic_po W=0.33 L=11 m=1
Rrespu2 PU_H_N int_res sky130_fd_pr__res_generic_po W=0.33 L=4 m=1
Xmnin_fast<3>_q0 net30 DRVHI_H int<3> net017<0> sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnin_fast<2>_q0 net30 DRVHI_H int<2> net017<1> sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnin_fast<1>_q0 net30 DRVHI_H int<1> net017<2> sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnin_fast<0>_q0 net30 DRVHI_H int<0> net017<3> sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnen_slow1_q0 n<2> PUEN_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=0.75 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnin_slow_q0 PU_H_N DRVHI_H n<2> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=0.42 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnen_fast<3>_q0 int<3> EN_FAST[3] VGND_IO net018<0>
+ sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xmnen_fast<2>_q0 int<2> EN_FAST[2] VGND_IO net018<1>
+ sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xmnen_fast<1>_q0 int<1> EN_FAST[1] VGND_IO net018<2>
+ sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xmnen_fast<0>_q0 int<0> EN_FAST[0] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5
+ m=1 w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpen_q0 PU_H_N PUEN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmpin_q0 PU_H_N DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=3 w=5.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_pupredrvr_strong_nd2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_ovtv2_pupredrvr_strong_nd3 DRVHI_H EN_FAST[3]
+ EN_FAST[2] EN_FAST[1] EN_FAST[0] PU_H_N PUEN_H VCC_IO VGND_IO
*.PININFO DRVHI_H:I EN_FAST[3]:I EN_FAST[2]:I EN_FAST[1]:I
*.PININFO EN_FAST[0]:I PU_H_N:O PUEN_H:I VCC_IO:I VGND_IO:I
XE1 net30 PU_H_N sky130_fd_io__tk_em1s
Rrespu1 int_res net30 sky130_fd_pr__res_generic_po W=0.33 L=11 m=1
Rrespu2 PU_H_N int_res sky130_fd_pr__res_generic_po W=0.33 L=4 m=1
Xmnin_fast<3>_q0 net30 DRVHI_H int<3> net017<0> sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnin_fast<2>_q0 net30 DRVHI_H int<2> net017<1> sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnin_fast<1>_q0 net30 DRVHI_H int<1> net017<2> sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnin_fast<0>_q0 net30 DRVHI_H int<0> net017<3> sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnen_slow1_q0 n<2> PUEN_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=0.75 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnin_slow_q0 PU_H_N DRVHI_H n<2> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=0.42 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnen_fast<3>_q0 int<3> EN_FAST[3] VGND_IO net018<0>
+ sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xmnen_fast<2>_q0 int<2> EN_FAST[2] VGND_IO net018<1>
+ sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xmnen_fast<1>_q0 int<1> EN_FAST[1] VGND_IO net018<2>
+ sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xmnen_fast<0>_q0 int<0> EN_FAST[0] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5
+ m=1 w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpen_q0 PU_H_N PUEN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmpin_q0 PU_H_N DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=3 w=5.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_ovtv2_pupredrvr_strong_nd3

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_pddrvr_strong FORCE_LO_H FORCE_LOVOL_H PAD PD_H[3]
+ PD_H[2] TIE_LO_ESD VCC_IO VGND_IO VSSIO_AMX
*.PININFO FORCE_LO_H:I FORCE_LOVOL_H:I PAD:O PD_H[3]:I PD_H[2]:I
*.PININFO TIE_LO_ESD:O VCC_IO:I VGND_IO:I VSSIO_AMX:I
XI112 PD_H[2] net61 sky130_fd_io__tk_em2s
XI113 PD_H[2] net59 sky130_fd_io__tk_em2s
XI97 PD_H[3] net85 sky130_fd_io__tk_em2s
XI108 TIE_LO_ESD net83 sky130_fd_io__tk_em2s
XI109 TIE_LO_ESD net77 sky130_fd_io__tk_em2s
XI102 PD_H[3] net73 sky130_fd_io__tk_em2s
XI104 PD_H[3] net69 sky130_fd_io__tk_em2s
XI96 PD_H[3] net67 sky130_fd_io__tk_em2s
XI87 TIE_LO_ESD net59 sky130_fd_io__tk_em2o
XI83 PD_H[3] net61 sky130_fd_io__tk_em2o
XI99 TIE_LO_ESD net85 sky130_fd_io__tk_em2o
XI82 TIE_LO_ESD net61 sky130_fd_io__tk_em2o
XI98 PD_H[2] net85 sky130_fd_io__tk_em2o
XI106 PD_H[2] net83 sky130_fd_io__tk_em2o
XI107 PD_H[3] net83 sky130_fd_io__tk_em2o
XI110 PD_H[3] net77 sky130_fd_io__tk_em2o
XI111 PD_H[2] net77 sky130_fd_io__tk_em2o
XI100 TIE_LO_ESD net73 sky130_fd_io__tk_em2o
XI101 PD_H[2] net73 sky130_fd_io__tk_em2o
XI103 TIE_LO_ESD net69 sky130_fd_io__tk_em2o
XI105 PD_H[2] net69 sky130_fd_io__tk_em2o
XI95 PD_H[2] net67 sky130_fd_io__tk_em2o
XI94 TIE_LO_ESD net67 sky130_fd_io__tk_em2o
XI88 PD_H[3] net59 sky130_fd_io__tk_em2o
XI49 VGND_IO TIE_LO_ESD sky130_fd_io__tk_tie_r_out_esd
Xn24<2>_q0 PAD net85 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn24<1>_q0 PAD net85 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn24<0>_q0 PAD net85 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn23<2>_q0 PAD net67 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn23<1>_q0 PAD net67 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn23<0>_q0 PAD net67 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn22<2>_q0 PAD PD_H[3] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn22<1>_q0 PAD PD_H[3] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn22<0>_q0 PAD PD_H[3] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn21<2>_q0 PAD PD_H[3] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn21<1>_q0 PAD PD_H[3] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn21<0>_q0 PAD PD_H[3] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn12_q0 PAD net61 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn32<2>_q0 PAD net69 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn32<1>_q0 PAD net69 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn32<0>_q0 PAD net69 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn33<2>_q0 PAD net83 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn33<1>_q0 PAD net83 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn33<0>_q0 PAD net83 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn34<3>_q0 PAD net77 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn34<2>_q0 PAD net77 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn34<1>_q0 PAD net77 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn34<0>_q0 PAD net77 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn11<2>_q0 PAD PD_H[2] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn11<1>_q0 PAD PD_H[2] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn11<0>_q0 PAD PD_H[2] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn13_q0 PAD net59 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn31_q0 PAD net73 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
xI72 VGND_IO VCC_IO sky130_fd_io__condiode
.ENDS sky130_fd_io__gpio_pddrvr_strong

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_pddrvr_strong_slow PAD PD_H VCC_IO VGND_IO
*.PININFO PAD:O PD_H:I VCC_IO:I VGND_IO:I
Xndrv_q0 PAD PD_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_pddrvr_strong_slow

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_pddrvr_weak PAD PD_H VCC_IO VGND_IO
*.PININFO PAD:O PD_H:I VCC_IO:I VGND_IO:I
Xndrv1_q0 PAD PD_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=6 w=5.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_pddrvr_weak

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_pudrvr_strong PAD PU_H_N[3] PU_H_N[2] TIE_HI_ESD
+ VCC_IO VNB
*.PININFO PAD:O PU_H_N[3]:I PU_H_N[2]:I TIE_HI_ESD:O VCC_IO:I VNB:I
XI112 PU_H_N[2] net43 sky130_fd_io__tk_em2s
XI108 TIE_HI_ESD net59 sky130_fd_io__tk_em2s
XI109 TIE_HI_ESD net53 sky130_fd_io__tk_em2s
XI104 PU_H_N[3] net49 sky130_fd_io__tk_em2s
XI125 PU_H_N[3] net45 sky130_fd_io__tk_em2s
XI83 PU_H_N[3] net43 sky130_fd_io__tk_em2o
XI82 TIE_HI_ESD net43 sky130_fd_io__tk_em2o
XI106 PU_H_N[2] net59 sky130_fd_io__tk_em2o
XI107 PU_H_N[3] net59 sky130_fd_io__tk_em2o
XI110 PU_H_N[3] net53 sky130_fd_io__tk_em2o
XI111 PU_H_N[2] net53 sky130_fd_io__tk_em2o
XI103 TIE_HI_ESD net49 sky130_fd_io__tk_em2o
XI105 PU_H_N[2] net49 sky130_fd_io__tk_em2o
XI124 TIE_HI_ESD net45 sky130_fd_io__tk_em2o
XI123 PU_H_N[2] net45 sky130_fd_io__tk_em2o
XI49 VCC_IO TIE_HI_ESD sky130_fd_io__tk_tie_r_out_esd
Xn24<2>_q0 PAD PU_H_N[3] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn24<1>_q0 PAD PU_H_N[3] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn24<0>_q0 PAD PU_H_N[3] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn23<2>_q0 PAD PU_H_N[3] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn23<1>_q0 PAD PU_H_N[3] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn23<0>_q0 PAD PU_H_N[3] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn22_q0 PAD net45 VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn21_q0 PAD PU_H_N[2] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn12<2>_q0 PAD net43 VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn12<1>_q0 PAD net43 VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn12<0>_q0 PAD net43 VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn32<2>_q0 PAD net49 VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn32<1>_q0 PAD net49 VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn32<0>_q0 PAD net49 VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn33<1>_q0 PAD net59 VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn33<0>_q0 PAD net59 VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn34<2>_q0 PAD net53 VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn34<1>_q0 PAD net53 VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn34<0>_q0 PAD net53 VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn11<2>_q0 PAD PU_H_N[2] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn11<1>_q0 PAD PU_H_N[2] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn11<0>_q0 PAD PU_H_N[2] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn13<2>_q0 PAD PU_H_N[2] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn13<1>_q0 PAD PU_H_N[2] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn13<0>_q0 PAD PU_H_N[2] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn31<2>_q0 PAD PU_H_N[3] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn31<1>_q0 PAD PU_H_N[3] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
Xn31<0>_q0 PAD PU_H_N[3] VCC_IO sky130_fd_io__gpio_pudrvr_unit_2_5
.ENDS sky130_fd_io__gpio_pudrvr_strong

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpio_pudrvr_unit_2_5 PD PGIN PS
*.PININFO PD:B PGIN:I PS:B
Xpdrv_q0 PD PGIN PS PS sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpio_pudrvr_unit_2_5

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux AMUXBUS_A AMUXBUS_B ANALOG_EN ANALOG_POL
+ ANALOG_SEL ENABLE_VDDA_H ENABLE_VSWITCH_H HLD_I_H HLD_I_H_N OUT PAD VCCD VDDA
+ VDDIO_Q VSSA VSSD VSSIO_Q VSWITCH
*.PININFO AMUXBUS_A:B AMUXBUS_B:B ANALOG_EN:I ANALOG_POL:I
*.PININFO ANALOG_SEL:I ENABLE_VDDA_H:I ENABLE_VSWITCH_H:I HLD_I_H:I
*.PININFO HLD_I_H_N:I OUT:I PAD:B VCCD:I VDDA:I VDDIO_Q:I VSSA:I
*.PININFO VSSD:I VSSIO_Q:I VSWITCH:I
xI43 VSSIO_Q VDDA sky130_fd_io__condiode
xI78 VSSA VSWITCH sky130_fd_io__condiode
Xmux_a_q0 AMUXBUS_A nga_amx_vpmp_h nga_pad_vpmp_h nmida_vccd net101 net101 net97
+ net97 net100 net99 net0127 HLD_I_H pga_amx_vdda_h_n pga_pad_vddioq_h_n VDDA
+ VDDIO_Q VSSA VSSD sky130_fd_io__gpiov2_amux_switch
Xmux_b_q0 AMUXBUS_B ngb_amx_vpmp_h ngb_pad_vpmp_h nmidb_vccd net101 net101 net97
+ net97 net100 net99 net0127 HLD_I_H pgb_amx_vdda_h_n pgb_pad_vddioq_h_n VDDA
+ VDDIO_Q VSSA VSSD sky130_fd_io__gpiov2_amux_switch
XBBM_logic ANALOG_EN ANALOG_POL ANALOG_SEL ENABLE_VDDA_H net0127
+ ENABLE_VSWITCH_H HLD_I_H HLD_I_H_N nga_amx_vpmp_h nga_pad_vpmp_h ngb_amx_vpmp_h
+ ngb_pad_vpmp_h nmida_vccd nmidb_vccd OUT pd_csd_vswitch_h pga_amx_vdda_h_n
+ pga_pad_vddioq_h_n pgb_amx_vdda_h_n pgb_pad_vddioq_h_n pu_csd_vddioq_h_n VCCD
+ VDDA VDDIO_Q VSSA VSSD VSWITCH sky130_fd_io__gpiov2_amux_ctl_logic
XI26 PAD net99 sky130_fd_io__res75only_small
XI58 net168 net97 sky130_fd_io__res75only_small
XI28 net166 net101 sky130_fd_io__res75only_small
XI57 PAD net168 sky130_fd_io__res75only_small
XI27 PAD net100 sky130_fd_io__res75only_small
XI55 PAD PAD sky130_fd_io__res75only_small
XI54 PAD net166 sky130_fd_io__res75only_small
XI53 PAD PAD sky130_fd_io__res75only_small
XI39 PAD net81 sky130_fd_io__res75only_small
XI40 PAD net85 sky130_fd_io__res75only_small
XI52 net81 pu_csd_vddioq_h_n VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=3
+ w=15.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XMP_PU net85 pu_csd_vddioq_h_n VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=4
+ w=15.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI49 net81 pd_csd_vswitch_h VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 m=6
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XMN_PD net85 pd_csd_vswitch_h VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 m=8
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
.ENDS sky130_fd_io__gpiov2_amux

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_ctl_inv_1 IN OUT VGND VPWR
*.PININFO IN:I OUT:O VGND:I VPWR:I
XI27 OUT IN VGND VGND sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI29 OUT IN VPWR VPWR sky130_fd_pr__pfet_01v8_hvt m=1 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amux_ctl_inv_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_ctl_logic ANALOG_EN ANALOG_POL ANALOG_SEL
+ ENABLE_VDDA_H ENABLE_VDDA_H_N ENABLE_VSWITCH_H HLD_I_H HLD_I_H_N
+ NGA_AMX_VSWITCH_H NGA_PAD_VSWITCH_H NGB_AMX_VSWITCH_H NGB_PAD_VSWITCH_H
+ NMIDA_VCCD NMIDB_VCCD OUT PD_CSD_VSWITCH_H PGA_AMX_VDDA_H_N PGA_PAD_VDDIOQ_H_N
+ PGB_AMX_VDDA_H_N PGB_PAD_VDDIOQ_H_N PU_CSD_VDDIOQ_H_N VCCD VDDA VDDIO_Q VSSA
+ VSSD VSWITCH
*.PININFO ANALOG_EN:I ANALOG_POL:I ANALOG_SEL:I ENABLE_VDDA_H:I
*.PININFO ENABLE_VDDA_H_N:O ENABLE_VSWITCH_H:I HLD_I_H:I HLD_I_H_N:I
*.PININFO NGA_AMX_VSWITCH_H:O NGA_PAD_VSWITCH_H:O NGB_AMX_VSWITCH_H:O
*.PININFO NGB_PAD_VSWITCH_H:O NMIDA_VCCD:O NMIDB_VCCD:O OUT:I
*.PININFO PD_CSD_VSWITCH_H:O PGA_AMX_VDDA_H_N:O PGA_PAD_VDDIOQ_H_N:O
*.PININFO PGB_AMX_VDDA_H_N:O PGB_PAD_VDDIOQ_H_N:O PU_CSD_VDDIOQ_H_N:O
*.PININFO VCCD:I VDDA:I VDDIO_Q:I VSSA:I VSSD:I VSWITCH:I
Xamux_sw_drvr_q0 amux_en_vdda_h amux_en_vdda_h_n amux_en_vddio_h
+ amux_en_vddio_h_n amux_en_vswitch_h amux_en_vswitch_h_n amuxbusa_on
+ amuxbusa_on_n amuxbusb_on amuxbusb_on_n NGA_AMX_VSWITCH_H NGA_PAD_VSWITCH_H
+ nga_pad_vswitch_h_n NGB_AMX_VSWITCH_H NGB_PAD_VSWITCH_H ngb_pad_vswitch_h_n
+ nmida_on_n NMIDA_VCCD nmida_vccd_n nmidb_on_n NMIDB_VCCD nmidb_vccd_n
+ PD_CSD_VSWITCH_H pd_csd_vswitch_h_n pd_on pd_on_n PGA_AMX_VDDA_H_N
+ PGA_PAD_VDDIOQ_H_N PGB_AMX_VDDA_H_N PGB_PAD_VDDIOQ_H_N PU_CSD_VDDIOQ_H_N pu_on
+ pu_on_n VCCD VDDA VDDIO_Q VSSA VSSD VSWITCH sky130_fd_io__gpiov2_amux_drvr
Xamux_lv_decoder_q0 amuxbusa_on amuxbusa_on_n amuxbusb_on amuxbusb_on_n
+ ANALOG_EN ANALOG_POL ANALOG_SEL NGA_PAD_VSWITCH_H nga_pad_vswitch_h_n
+ NGB_PAD_VSWITCH_H ngb_pad_vswitch_h_n nmida_on_n nmida_vccd_n nmidb_on_n
+ nmidb_vccd_n OUT pd_on pd_on_n pd_csd_vswitch_h_n PGA_AMX_VDDA_H_N
+ PGA_PAD_VDDIOQ_H_N PGB_AMX_VDDA_H_N PGB_PAD_VDDIOQ_H_N pu_on pu_on_n
+ PU_CSD_VDDIOQ_H_N VCCD VSSD sky130_fd_io__gpiov2_amux_decoder
Xamux_ls_q0 amux_en_vdda_h amux_en_vdda_h_n amux_en_vddio_h amux_en_vddio_h_n
+ amux_en_vswitch_h amux_en_vswitch_h_n ANALOG_EN ENABLE_VDDA_H ENABLE_VDDA_H_N
+ ENABLE_VSWITCH_H HLD_I_H HLD_I_H_N VCCD VDDA VDDIO_Q VSSA VSSD VSWITCH
+ sky130_fd_io__gpiov2_amux_ls
.ENDS sky130_fd_io__gpiov2_amux_ctl_logic

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_ctl_logic_i2c_fix ANALOG_EN ANALOG_POL
+ ANALOG_SEL ENABLE_VDDA_H ENABLE_VDDA_H_N ENABLE_VSWITCH_H HLD_I_H_N
+ NGA_AMX_VSWITCH_H NGA_PAD_VSWITCH_H NGB_AMX_VSWITCH_H NGB_PAD_VSWITCH_H
+ NMIDA_VCCD NMIDB_VCCD OUT PD_CSD_VSWITCH_H PGA_AMX_VDDA_H_N PGA_PAD_VDDIOQ_H_N
+ PGB_AMX_VDDA_H_N PGB_PAD_VDDIOQ_H_N PU_CSD_VDDIOQ_H_N VCCD VDDA VDDIO_Q VSSA
+ VSSD VSWITCH
*.PININFO ANALOG_EN:I ANALOG_POL:I ANALOG_SEL:I ENABLE_VDDA_H:I
*.PININFO ENABLE_VDDA_H_N:O ENABLE_VSWITCH_H:I HLD_I_H_N:I
*.PININFO NGA_AMX_VSWITCH_H:O NGA_PAD_VSWITCH_H:O NGB_AMX_VSWITCH_H:O
*.PININFO NGB_PAD_VSWITCH_H:O NMIDA_VCCD:O NMIDB_VCCD:O OUT:I
*.PININFO PD_CSD_VSWITCH_H:O PGA_AMX_VDDA_H_N:O PGA_PAD_VDDIOQ_H_N:O
*.PININFO PGB_AMX_VDDA_H_N:O PGB_PAD_VDDIOQ_H_N:O PU_CSD_VDDIOQ_H_N:O
*.PININFO VCCD:I VDDA:I VDDIO_Q:I VSSA:I VSSD:I VSWITCH:I
Xamux_ls_q0 amux_en_vdda_h amux_en_vdda_h_n amux_en_vddio_h amux_en_vswitch_h
+ amux_en_vswitch_h_n ANALOG_EN ENABLE_VDDA_H ENABLE_VDDA_H_N ENABLE_VSWITCH_H
+ HLD_I_H_N VCCD VDDA VDDIO_Q VSSA VSSD VSWITCH
+ sky130_fd_io__gpiov2_amux_ls_i2c_fix
Xamux_sw_drvr_q0 amux_en_vdda_h amux_en_vdda_h_n amux_en_vddio_h
+ amux_en_vswitch_h amux_en_vswitch_h_n amuxbusa_on amuxbusa_on_n amuxbusb_on
+ amuxbusb_on_n HLD_I_H_N NGA_AMX_VSWITCH_H NGA_PAD_VSWITCH_H nga_pad_vswitch_h_n
+ NGB_AMX_VSWITCH_H NGB_PAD_VSWITCH_H ngb_pad_vswitch_h_n nmida_on_n NMIDA_VCCD
+ nmida_vccd_n nmidb_on_n NMIDB_VCCD nmidb_vccd_n PD_CSD_VSWITCH_H
+ pd_csd_vswitch_h_n pd_on pd_on_n PGA_AMX_VDDA_H_N PGA_PAD_VDDIOQ_H_N
+ PGB_AMX_VDDA_H_N PGB_PAD_VDDIOQ_H_N PU_CSD_VDDIOQ_H_N pu_on pu_on_n VCCD VDDA
+ VDDIO_Q VSSA VSSD VSWITCH sky130_fd_io__gpiov2_amux_drvr_i2c_fix
Xamux_lv_decoder_q0 amuxbusa_on amuxbusa_on_n amuxbusb_on amuxbusb_on_n
+ ANALOG_EN ANALOG_POL ANALOG_SEL NGA_PAD_VSWITCH_H nga_pad_vswitch_h_n
+ NGB_PAD_VSWITCH_H ngb_pad_vswitch_h_n nmida_on_n nmida_vccd_n nmidb_on_n
+ nmidb_vccd_n OUT pd_on pd_on_n pd_csd_vswitch_h_n PGA_AMX_VDDA_H_N
+ PGA_PAD_VDDIOQ_H_N PGB_AMX_VDDA_H_N PGB_PAD_VDDIOQ_H_N pu_on pu_on_n
+ PU_CSD_VDDIOQ_H_N VCCD VSSD sky130_fd_io__gpiov2_amux_decoder
.ENDS sky130_fd_io__gpiov2_amux_ctl_logic_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_ctl_ls IN IN_B OUT_H OUT_H_N RST_H RST_H_N
+ VGND VPWR_HV VPWR_LV
*.PININFO IN:I IN_B:I OUT_H:O OUT_H_N:O RST_H:I RST_H_N:I VGND:I
*.PININFO VPWR_HV:I VPWR_LV:I
XI14 OUT_H fbk_n VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI11 OUT_H_N fbk VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 fbk_n fbk VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 fbk fbk_n VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI5 net61 RST_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=4 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI13 OUT_H fbk_n VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 OUT_H_N fbk VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI58 fbk VPWR_LV net62 VGND sky130_fd_pr__nfet_05v0_nvt m=4 w=1.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmnrst_q0 fbk RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI59 fbk_n VPWR_LV net66 VGND sky130_fd_pr__nfet_05v0_nvt m=4 w=1.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI8 net66 IN net61 VGND sky130_fd_pr__nfet_01v8_lvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI7 net62 IN_B net61 VGND sky130_fd_pr__nfet_01v8_lvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amux_ctl_ls

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_ctl_ls_i2c_fix IN IN_B OUT_H RST_H RST_H_N
+ VGND VPWR_HV VPWR_LV
*.PININFO IN:I IN_B:I OUT_H:O RST_H:I RST_H_N:I VGND:I VPWR_HV:I
*.PININFO VPWR_LV:I
XI14 fbk_n RST_H_N VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=2 w=0.75 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI11 OUT_H fbk_n VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=2 w=0.75 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 fbk_n fbk VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 fbk fbk_n VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI5 net70 RST_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=4 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 OUT_H fbk_n VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI58 fbk VPWR_LV net71 VGND sky130_fd_pr__nfet_05v0_nvt m=4 w=1.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmnrst_q0 fbk RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI59 fbk_n VPWR_LV net75 VGND sky130_fd_pr__nfet_05v0_nvt m=4 w=1.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI8 net75 IN net70 VGND sky130_fd_pr__nfet_01v8_lvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI7 net71 IN_B net70 VGND sky130_fd_pr__nfet_01v8_lvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amux_ctl_ls_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_ctl_lshv2hv IN IN_B OUT_H OUT_H_N RST_H
+ RST_H_N VGND VPWR_HV
*.PININFO IN:I IN_B:I OUT_H:O OUT_H_N:O RST_H:I RST_H_N:I VGND:I
*.PININFO VPWR_HV:I
XI14 OUT_H_N fbk VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI11 OUT_H fbk_n VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 fbk fbk_n VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 fbk_n fbk VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI64 net64 RST_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI13 OUT_H_N fbk VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 OUT_H fbk_n VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmnrst_q0 fbk RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI8 fbk_n IN net64 VGND sky130_fd_pr__nfet_g5v0d10v5 m=3 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI7 fbk IN_B net64 VGND sky130_fd_pr__nfet_g5v0d10v5 m=3 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amux_ctl_lshv2hv

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_decoder AMUXBUSA_ON AMUXBUSA_ON_N AMUXBUSB_ON
+ AMUXBUSB_ON_N ANALOG_EN ANALOG_POL ANALOG_SEL NGA_PAD_VSWITCH_H
+ NGA_PAD_VSWITCH_H_N NGB_PAD_VSWITCH_H NGB_PAD_VSWITCH_H_N NMIDA_ON_N
+ NMIDA_VCCD_N D_B NMIDB_VCCD_N OUT PD_ON PD_ON_N PD_VSWITCH_H_N PGA_AMX_VDDA_H_N
+ PGA_PAD_VDDIOQ_H_N PGB_AMX_VDDA_H_N PGB_PAD_VDDIOQ_H_N PU_ON PU_ON_N
+ PU_VDDIOQ_H_N VCCD VSSD
*.PININFO AMUXBUSA_ON:O AMUXBUSA_ON_N:O AMUXBUSB_ON:O AMUXBUSB_ON_N:O
*.PININFO ANALOG_EN:I ANALOG_POL:I ANALOG_SEL:I NGA_PAD_VSWITCH_H:I
*.PININFO NGA_PAD_VSWITCH_H_N:I NGB_PAD_VSWITCH_H:I
*.PININFO NGB_PAD_VSWITCH_H_N:I NMIDA_ON_N:O NMIDA_VCCD_N:I D_B:O
*.PININFO NMIDB_VCCD_N:I OUT:I PD_ON:O PD_ON_N:O PD_VSWITCH_H_N:I
*.PININFO PGA_AMX_VDDA_H_N:I PGA_PAD_VDDIOQ_H_N:I PGB_AMX_VDDA_H_N:I
*.PININFO PGB_PAD_VDDIOQ_H_N:I PU_ON:O PU_ON_N:O PU_VDDIOQ_H_N:I
*.PININFO VCCD:I VSSD:I
XI116 ana_en_i_n int_pd_on_n int_pd_on VSSD VSSD VCCD VCCD sky130_fd_io__nor2_1
XI113 ana_en_i_n net144 int_amuxa_on VSSD VSSD VCCD VCCD sky130_fd_io__nor2_1
XI115 ana_en_i_n int_pu_on_n int_pu_on VSSD VSSD VCCD VCCD sky130_fd_io__nor2_1
XI114 ana_en_i_n net137 int_amuxb_on VSSD VSSD VCCD VCCD sky130_fd_io__nor2_1
XI111 ana_pol_i out_i int_pu_on_n VSSD VSSD VCCD VCCD sky130_fd_io__nand2_1
XI112 ana_pol_i_n out_i_n int_pd_on_n VSSD VSSD VCCD VCCD sky130_fd_io__nand2_1
XI109 ana_sel_i_n pol_xor_out net144 VSSD VSSD VCCD VCCD sky130_fd_io__nand2_1
XI110 pol_xor_out ana_sel_i net137 VSSD VSSD VCCD VCCD sky130_fd_io__nand2_1
XI106 NGB_PAD_VSWITCH_H net212 net172 VSSD VCCD sky130_fd_io__hvsbt_nor
XI102 NGA_PAD_VSWITCH_H net222 net167 VSSD VCCD sky130_fd_io__hvsbt_nor
XI79 int_pu_on PGA_PAD_VDDIOQ_H_N PGB_PAD_VDDIOQ_H_N NGA_PAD_VSWITCH_H_N
+ NGB_PAD_VSWITCH_H_N int_fbk_puon_n VSSD VCCD sky130_fd_io__gpiov2_amux_nand5
XI80 int_pd_on PGA_PAD_VDDIOQ_H_N PGB_PAD_VDDIOQ_H_N NGA_PAD_VSWITCH_H_N
+ NGB_PAD_VSWITCH_H_N int_fbk_pdon_n VSSD VCCD sky130_fd_io__gpiov2_amux_nand5
XI78 int_amuxb_on PU_VDDIOQ_H_N PD_VSWITCH_H_N NMIDB_VCCD_N AMUXBUSB_ON_N VSSD
+ VCCD sky130_fd_io__gpiov2_amux_nand4
XI77 int_amuxa_on PU_VDDIOQ_H_N PD_VSWITCH_H_N NMIDA_VCCD_N AMUXBUSA_ON_N VSSD
+ VCCD sky130_fd_io__gpiov2_amux_nand4
XI101 PGA_PAD_VDDIOQ_H_N PGA_AMX_VDDA_H_N net222 VSSD VCCD
+ sky130_fd_io__hvsbt_nand2
XI121 int_amux_b_on_n net172 D_B VSSD VCCD sky130_fd_io__hvsbt_nand2
XI105 PGB_PAD_VDDIOQ_H_N PGB_AMX_VDDA_H_N net212 VSSD VCCD
+ sky130_fd_io__hvsbt_nand2
XI120 int_amux_a_on_n net167 NMIDA_ON_N VSSD VCCD sky130_fd_io__hvsbt_nand2
XI45 ana_pol_i out_i pol_xor_out VSSD VCCD sky130_fd_io__xor2_1
XI41 ana_pol_i_n ana_pol_i VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
XI89 int_amuxa_on int_amux_a_on_n VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
XI39 ANALOG_SEL ana_sel_i_n VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
XI40 ana_sel_i_n ana_sel_i VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
XI35 ANALOG_POL ana_pol_i_n VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
XI74 AMUXBUSB_ON_N AMUXBUSB_ON VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
XI73 AMUXBUSA_ON_N AMUXBUSA_ON VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
XI76 int_fbk_pdon_n PD_ON VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
XI58 ANALOG_EN ana_en_i_n VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
XI75 int_fbk_puon_n PU_ON VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
XI43 OUT out_i_n VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
XI44 out_i_n out_i VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
XI91 int_amuxb_on int_amux_b_on_n VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
XI93 PU_ON PU_ON_N VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
XI95 PD_ON PD_ON_N VSSD VSSD VCCD VCCD sky130_fd_io__inv_1
.ENDS sky130_fd_io__gpiov2_amux_decoder

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_drvr AMUX_EN_VDDA_H AMUX_EN_VDDA_H_N
+ AMUX_EN_VDDIO_H AMUX_EN_VDDIO_H_N AMUX_EN_VSWITCH_H AMUX_EN_VSWITCH_H_N
+ AMUXBUSA_ON AMUXBUSA_ON_N AMUXBUSB_ON AMUXBUSB_ON_N NGA_AMX_VSWITCH_H
+ NGA_PAD_VSWITCH_H NGA_PAD_VSWITCH_H_N NGB_AMX_VSWITCH_H NGB_PAD_VSWITCH_H
+ NGB_PAD_VSWITCH_H_N NMIDA_ON_N NMIDA_VCCD NMIDA_VCCD_N D_B NMIDB_VCCD
+ NMIDB_VCCD_N PD_CSD_VSWITCH_H PD_CSD_VSWITCH_H_N PD_ON PD_ON_N PGA_AMX_VDDA_H_N
+ PGA_PAD_VDDIOQ_H_N PGB_AMX_VDDA_H_N PGB_PAD_VDDIOQ_H_N PU_CSD_VDDIOQ_H_N PU_ON
+ PU_ON_N VCCD VDDA VDDIO_Q VSSA VSSD VSWITCH
*.PININFO AMUX_EN_VDDA_H:I AMUX_EN_VDDA_H_N:I AMUX_EN_VDDIO_H:I
*.PININFO AMUX_EN_VDDIO_H_N:I AMUX_EN_VSWITCH_H:I
*.PININFO AMUX_EN_VSWITCH_H_N:I AMUXBUSA_ON:I AMUXBUSA_ON_N:I
*.PININFO AMUXBUSB_ON:I AMUXBUSB_ON_N:I NGA_AMX_VSWITCH_H:O
*.PININFO NGA_PAD_VSWITCH_H:O NGA_PAD_VSWITCH_H_N:O
*.PININFO NGB_AMX_VSWITCH_H:O NGB_PAD_VSWITCH_H:O
*.PININFO NGB_PAD_VSWITCH_H_N:O NMIDA_ON_N:I NMIDA_VCCD:O
*.PININFO NMIDA_VCCD_N:O D_B:I NMIDB_VCCD:O NMIDB_VCCD_N:O
*.PININFO PD_CSD_VSWITCH_H:O PD_CSD_VSWITCH_H_N:O PD_ON:I PD_ON_N:I
*.PININFO PGA_AMX_VDDA_H_N:O PGA_PAD_VDDIOQ_H_N:O PGB_AMX_VDDA_H_N:O
*.PININFO PGB_PAD_VDDIOQ_H_N:O PU_CSD_VDDIOQ_H_N:O PU_ON:I PU_ON_N:I
*.PININFO VCCD:I VDDA:I VDDIO_Q:I VSSA:I VSSD:I VSWITCH:I
XI93 NMIDA_VCCD NMIDA_VCCD_N VSSD VCCD sky130_fd_io__hvsbt_inv_x1
XI105 NMIDB_VCCD NMIDB_VCCD_N VSSD VCCD sky130_fd_io__hvsbt_inv_x1
XI38 net274 PU_CSD_VDDIOQ_H_N VDDIO_Q VSSD sky130_fd_io__gpiov2_amx_pucsd_inv
Xpga_amx_ls_q0 net265 net272 PGA_AMX_VDDA_H_N AMUX_EN_VDDA_H_N AMUX_EN_VDDA_H
+ VSSA VDDA sky130_fd_io__gpiov2_amux_drvr_lshv2hv
XI103 net239 net245 PGB_AMX_VDDA_H_N AMUX_EN_VDDA_H_N AMUX_EN_VDDA_H VSSA VDDA
+ sky130_fd_io__gpiov2_amux_drvr_lshv2hv
XI45 net256 NGA_AMX_VSWITCH_H VSWITCH VSSA sky130_fd_io__gpiov2_amx_inv4
XI42 net265 PGA_PAD_VDDIOQ_H_N VDDIO_Q VSSD sky130_fd_io__gpiov2_amx_inv4
XI47 net256 NGA_PAD_VSWITCH_H VSWITCH VSSA sky130_fd_io__gpiov2_amx_inv4
XI62 net239 PGB_PAD_VDDIOQ_H_N VDDIO_Q VSSD sky130_fd_io__gpiov2_amx_inv4
XI63 net236 NGB_AMX_VSWITCH_H VSWITCH VSSA sky130_fd_io__gpiov2_amx_inv4
XI64 net236 NGB_PAD_VSWITCH_H VSWITCH VSSA sky130_fd_io__gpiov2_amx_inv4
XI53 D_B NMIDB_VCCD VSSD VCCD sky130_fd_io__hvsbt_inv_x2
XI89 NMIDA_ON_N NMIDA_VCCD VSSD VCCD sky130_fd_io__hvsbt_inv_x2
Xpdcsd_inv_q0 net254 PD_CSD_VSWITCH_H VSWITCH VSSA
+ sky130_fd_io__gpiov2_amx_pdcsd_inv
XI90 PD_CSD_VSWITCH_H PD_CSD_VSWITCH_H_N VSWITCH VSSA sky130_fd_io__amx_inv1
XI85 NGB_PAD_VSWITCH_H NGB_PAD_VSWITCH_H_N VSWITCH VSSA sky130_fd_io__amx_inv1
XI87 NGA_PAD_VSWITCH_H NGA_PAD_VSWITCH_H_N VSWITCH VSSA sky130_fd_io__amx_inv1
Xpu_csd_ls_q0 PU_ON PU_ON_N net274 net275 AMUX_EN_VDDIO_H_N AMUX_EN_VDDIO_H VSSD
+ VDDIO_Q VCCD sky130_fd_io__gpiov2_amux_drvr_ls
Xpga_pad_ls_q0 AMUXBUSA_ON AMUXBUSA_ON_N net265 net272 AMUX_EN_VDDIO_H_N
+ AMUX_EN_VDDIO_H VSSD VDDIO_Q VCCD sky130_fd_io__gpiov2_amux_drvr_ls
Xnga_ls_q0 AMUXBUSA_ON AMUXBUSA_ON_N net257 net256 AMUX_EN_VSWITCH_H_N
+ AMUX_EN_VSWITCH_H VSSA VSWITCH VCCD sky130_fd_io__gpiov2_amux_drvr_ls
Xpd_csd_ls_q0 PD_ON PD_ON_N net248 net254 AMUX_EN_VSWITCH_H_N AMUX_EN_VSWITCH_H
+ VSSA VSWITCH VCCD sky130_fd_io__gpiov2_amux_drvr_ls
Xpgb_pad_ls_q0 AMUXBUSB_ON AMUXBUSB_ON_N net239 net245 AMUX_EN_VDDIO_H_N
+ AMUX_EN_VDDIO_H VSSD VDDIO_Q VCCD sky130_fd_io__gpiov2_amux_drvr_ls
Xngb_ls_q0 AMUXBUSB_ON AMUXBUSB_ON_N net230 net236 AMUX_EN_VSWITCH_H_N
+ AMUX_EN_VSWITCH_H VSSA VSWITCH VCCD sky130_fd_io__gpiov2_amux_drvr_ls
XI76 NGB_AMX_VSWITCH_H AMUX_EN_VDDA_H_N VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5
+ m=1 w=1.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI77 NGB_PAD_VSWITCH_H AMUX_EN_VDDIO_H_N VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5
+ m=1 w=1.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI75 NGA_AMX_VSWITCH_H AMUX_EN_VDDA_H_N VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5
+ m=1 w=1.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI78 NGA_PAD_VSWITCH_H AMUX_EN_VDDIO_H_N VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5
+ m=1 w=1.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI104 PD_CSD_VSWITCH_H AMUX_EN_VDDIO_H_N VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5
+ m=1 w=1.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
.ENDS sky130_fd_io__gpiov2_amux_drvr

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_drvr_i2c_fix AMUX_EN_VDDA_H AMUX_EN_VDDA_H_N
+ AMUX_EN_VDDIO_H AMUX_EN_VSWITCH_H AMUX_EN_VSWITCH_H_N AMUXBUSA_ON AMUXBUSA_ON_N
+ AMUXBUSB_ON AMUXBUSB_ON_N HLD_I_H_N NGA_AMX_VSWITCH_H NGA_PAD_VSWITCH_H
+ NGA_PAD_VSWITCH_H_N NGB_AMX_VSWITCH_H NGB_PAD_VSWITCH_H NGB_PAD_VSWITCH_H_N
+ NMIDA_ON_N NMIDA_VCCD NMIDA_VCCD_N D_B NMIDB_VCCD NMIDB_VCCD_N PD_CSD_VSWITCH_H
+ PD_CSD_VSWITCH_H_N PD_ON PD_ON_N PGA_AMX_VDDA_H_N PGA_PAD_VDDIOQ_H_N
+ PGB_AMX_VDDA_H_N PGB_PAD_VDDIOQ_H_N PU_CSD_VDDIOQ_H_N PU_ON PU_ON_N VCCD VDDA
+ VDDIO_Q VSSA VSSD VSWITCH
*.PININFO AMUX_EN_VDDA_H:I AMUX_EN_VDDA_H_N:I AMUX_EN_VDDIO_H:I
*.PININFO AMUX_EN_VSWITCH_H:I AMUX_EN_VSWITCH_H_N:I AMUXBUSA_ON:I
*.PININFO AMUXBUSA_ON_N:I AMUXBUSB_ON:I AMUXBUSB_ON_N:I HLD_I_H_N:I
*.PININFO NGA_AMX_VSWITCH_H:O NGA_PAD_VSWITCH_H:O
*.PININFO NGA_PAD_VSWITCH_H_N:O NGB_AMX_VSWITCH_H:O
*.PININFO NGB_PAD_VSWITCH_H:O NGB_PAD_VSWITCH_H_N:O NMIDA_ON_N:I
*.PININFO NMIDA_VCCD:O NMIDA_VCCD_N:O D_B:I NMIDB_VCCD:O
*.PININFO NMIDB_VCCD_N:O PD_CSD_VSWITCH_H:O PD_CSD_VSWITCH_H_N:O
*.PININFO PD_ON:I PD_ON_N:I PGA_AMX_VDDA_H_N:O PGA_PAD_VDDIOQ_H_N:O
*.PININFO PGB_AMX_VDDA_H_N:O PGB_PAD_VDDIOQ_H_N:O PU_CSD_VDDIOQ_H_N:O
*.PININFO PU_ON:I PU_ON_N:I VCCD:I VDDA:I VDDIO_Q:I VSSA:I VSSD:I
*.PININFO VSWITCH:I
Xpga_pad_ls_q0 AMUXBUSA_ON AMUXBUSA_ON_N net154 net160 hld_i_h HLD_I_H_N
+ amux_en_vddio_h_n AMUX_EN_VDDIO_H VSSD VDDIO_Q VCCD
+ sky130_fd_io__gpiov2_amux_drvr_ls_i2c_fix3_ver2
Xpgb_pad_ls_q0 AMUXBUSB_ON AMUXBUSB_ON_N net144 net149 hld_i_h HLD_I_H_N
+ amux_en_vddio_h_n AMUX_EN_VDDIO_H VSSD VDDIO_Q VCCD
+ sky130_fd_io__gpiov2_amux_drvr_ls_i2c_fix3_ver2
XI38 net168 PU_CSD_VDDIOQ_H_N VDDIO_Q VSSD sky130_fd_io__gpiov2_amx_pucsd_buf
Xpu_csd_ls_q0 PU_ON PU_ON_N net167 net168 HLD_I_H_N AMUX_EN_VDDIO_H VSSD VDDIO_Q
+ VCCD sky130_fd_io__gpiov2_amux_drvr_ls_i2c_fix3
XI111 HLD_I_H_N hld_i_h VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
XI110 AMUX_EN_VDDIO_H amux_en_vddio_h_n VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
XI93 NMIDA_VCCD NMIDA_VCCD_N VSSD VCCD sky130_fd_io__hvsbt_inv_x1
XI105 NMIDB_VCCD NMIDB_VCCD_N VSSD VCCD sky130_fd_io__hvsbt_inv_x1
Xpga_amx_ls_q0 net154 net160 PGA_AMX_VDDA_H_N AMUX_EN_VDDA_H_N AMUX_EN_VDDA_H
+ VSSA VDDA sky130_fd_io__gpiov2_amux_drvr_lshv2hv
XI103 net144 net149 PGB_AMX_VDDA_H_N AMUX_EN_VDDA_H_N AMUX_EN_VDDA_H VSSA VDDA
+ sky130_fd_io__gpiov2_amux_drvr_lshv2hv
XI45 net295 NGA_AMX_VSWITCH_H VSWITCH VSSA sky130_fd_io__gpiov2_amx_inv4
XI42 net154 PGA_PAD_VDDIOQ_H_N VDDIO_Q VSSD sky130_fd_io__gpiov2_amx_inv4
XI47 net295 NGA_PAD_VSWITCH_H VSWITCH VSSA sky130_fd_io__gpiov2_amx_inv4
XI62 net144 PGB_PAD_VDDIOQ_H_N VDDIO_Q VSSD sky130_fd_io__gpiov2_amx_inv4
XI63 net284 NGB_AMX_VSWITCH_H VSWITCH VSSA sky130_fd_io__gpiov2_amx_inv4
XI64 net284 NGB_PAD_VSWITCH_H VSWITCH VSSA sky130_fd_io__gpiov2_amx_inv4
XI53 D_B NMIDB_VCCD VSSD VCCD sky130_fd_io__hvsbt_inv_x2
XI89 NMIDA_ON_N NMIDA_VCCD VSSD VCCD sky130_fd_io__hvsbt_inv_x2
Xpdcsd_inv_q0 net293 PD_CSD_VSWITCH_H VSWITCH VSSA
+ sky130_fd_io__gpiov2_amx_pdcsd_inv
XI87 NGA_PAD_VSWITCH_H NGA_PAD_VSWITCH_H_N VSWITCH VSSA sky130_fd_io__amx_inv1
XI85 NGB_PAD_VSWITCH_H NGB_PAD_VSWITCH_H_N VSWITCH VSSA sky130_fd_io__amx_inv1
XI90 PD_CSD_VSWITCH_H PD_CSD_VSWITCH_H_N VSWITCH VSSA sky130_fd_io__amx_inv1
Xnga_ls_q0 AMUXBUSA_ON AMUXBUSA_ON_N net296 net295 AMUX_EN_VSWITCH_H_N
+ AMUX_EN_VSWITCH_H VSSA VSWITCH VCCD sky130_fd_io__gpiov2_amux_drvr_ls
Xpd_csd_ls_q0 PD_ON PD_ON_N net287 net293 AMUX_EN_VSWITCH_H_N AMUX_EN_VSWITCH_H
+ VSSA VSWITCH VCCD sky130_fd_io__gpiov2_amux_drvr_ls
Xngb_ls_q0 AMUXBUSB_ON AMUXBUSB_ON_N net278 net284 AMUX_EN_VSWITCH_H_N
+ AMUX_EN_VSWITCH_H VSSA VSWITCH VCCD sky130_fd_io__gpiov2_amux_drvr_ls
XI76 NGB_AMX_VSWITCH_H AMUX_EN_VDDA_H_N VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5
+ m=1 w=1.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI77 NGB_PAD_VSWITCH_H amux_en_vddio_h_n VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5
+ m=1 w=1.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI75 NGA_AMX_VSWITCH_H AMUX_EN_VDDA_H_N VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5
+ m=1 w=1.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI78 NGA_PAD_VSWITCH_H amux_en_vddio_h_n VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5
+ m=1 w=1.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI104 PD_CSD_VSWITCH_H amux_en_vddio_h_n VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5
+ m=1 w=1.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
.ENDS sky130_fd_io__gpiov2_amux_drvr_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_drvr_ls IN IN_B OUT_H OUT_H_N RST_H RST_H_N
+ VGND VPWR_HV VPWR_LV
*.PININFO IN:I IN_B:I OUT_H:O OUT_H_N:O RST_H:I RST_H_N:I VGND:I
*.PININFO VPWR_HV:I VPWR_LV:I
XI11 OUT_H_N OUT_H VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.7 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI9 OUT_H OUT_H_N VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.7 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI21 net42 VPWR_LV net58 VGND sky130_fd_pr__nfet_05v0_nvt m=2 w=1.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI20 net38 VPWR_LV net54 VGND sky130_fd_pr__nfet_05v0_nvt m=2 w=1.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI17 OUT_H RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.5 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 net58 IN VGND VGND sky130_fd_pr__nfet_01v8_lvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 net54 IN_B VGND VGND sky130_fd_pr__nfet_01v8_lvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI25 OUT_H RST_H_N net38 VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI24 OUT_H_N RST_H_N net42 VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amux_drvr_ls

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_drvr_ls_i2c_fix3 IN IN_B OUT_H OUT_H_N
+ RST2_H_N RST_H_N VGND VPWR_HV VPWR_LV
*.PININFO IN:I IN_B:I OUT_H:O OUT_H_N:O RST2_H_N:I RST_H_N:I VGND:I
*.PININFO VPWR_HV:I VPWR_LV:I
XI34 RST_H_N net086 VGND VPWR_HV sky130_fd_io__hvsbt_inv_x1
XI33 RST2_H_N net074 VGND VPWR_HV sky130_fd_io__hvsbt_inv_x1
XI11 OUT_H_N OUT_H VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.7 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI9 OUT_H OUT_H_N VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.7 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI29 OUT_H_N RST2_H_N VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=3 w=1.5
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI28 OUT_H_N RST_H_N VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI21 net55 VPWR_LV net79 VGND sky130_fd_pr__nfet_05v0_nvt m=2 w=1.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI20 net51 VPWR_LV net75 VGND sky130_fd_pr__nfet_05v0_nvt m=2 w=1.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI17 OUT_H net086 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 net79 IN VGND VGND sky130_fd_pr__nfet_01v8_lvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 net75 IN_B VGND VGND sky130_fd_pr__nfet_01v8_lvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI31 OUT_H net074 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.5 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI25 OUT_H RST_H_N net51 VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI24 OUT_H_N RST_H_N net55 VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amux_drvr_ls_i2c_fix3

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_drvr_ls_i2c_fix3_ver2 IN IN_B OUT_H OUT_H_N
+ RST2_H RST2_H_N RST_H RST_H_N VGND VPWR_HV VPWR_LV
*.PININFO IN:I IN_B:I OUT_H:O OUT_H_N:O RST2_H:I RST2_H_N:I RST_H:I
*.PININFO RST_H_N:I VGND:I VPWR_HV:I VPWR_LV:I
XI11 OUT_H_N OUT_H VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.7 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI9 OUT_H OUT_H_N VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.7 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI29 OUT_H_N RST2_H_N VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=3 w=1.5
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI28 OUT_H_N RST_H_N VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI21 net56 VPWR_LV net76 VGND sky130_fd_pr__nfet_05v0_nvt m=2 w=1.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI20 net52 VPWR_LV net72 VGND sky130_fd_pr__nfet_05v0_nvt m=2 w=1.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI17 OUT_H RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 net76 IN VGND VGND sky130_fd_pr__nfet_01v8_lvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 net72 IN_B VGND VGND sky130_fd_pr__nfet_01v8_lvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI31 OUT_H RST2_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.5 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI25 OUT_H RST_H_N net52 VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI24 OUT_H_N RST_H_N net56 VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amux_drvr_ls_i2c_fix3_ver2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_drvr_lshv2hv IN IN_B OUT_H_N RST_H RST_H_N
+ VGND VPWR_HV
*.PININFO IN:I IN_B:I OUT_H_N:O RST_H:I RST_H_N:I VGND:I VPWR_HV:I
XI14 OUT_H_N fbk VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 fbk fbk_n VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 fbk_n fbk VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI64 net52 RST_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI13 OUT_H_N fbk VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmnrst_q0 fbk RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI8 fbk_n IN net52 VGND sky130_fd_pr__nfet_g5v0d10v5 m=3 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI7 fbk IN_B net52 VGND sky130_fd_pr__nfet_g5v0d10v5 m=3 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amux_drvr_lshv2hv

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_ls AMUX_EN_VDDA_H AMUX_EN_VDDA_H_N
+ AMUX_EN_VDDIO_H AMUX_EN_VDDIO_H_N AMUX_EN_VSWITCH_H AMUX_EN_VSWITCH_H_N
+ ANALOG_EN ENABLE_VDDA_H ENABLE_VDDA_H_N ENABLE_VSWITCH_H HLD_I_H HLD_I_H_N VCCD
+ VDDA VDDIO_Q VSSA VSSD VSWITCH
*.PININFO AMUX_EN_VDDA_H:O AMUX_EN_VDDA_H_N:O AMUX_EN_VDDIO_H:O
*.PININFO AMUX_EN_VDDIO_H_N:O AMUX_EN_VSWITCH_H:O
*.PININFO AMUX_EN_VSWITCH_H_N:O ANALOG_EN:I ENABLE_VDDA_H:I
*.PININFO ENABLE_VDDA_H_N:O ENABLE_VSWITCH_H:I HLD_I_H:I HLD_I_H_N:I
*.PININFO VCCD:I VDDA:I VDDIO_Q:I VSSA:I VSSD:I VSWITCH:I
XI32 ENABLE_VDDA_H ENABLE_VDDA_H_N VSSA VDDA sky130_fd_io__gpiov2_amux_ls_inv_x1
Xpd_vswitch_ls_q0 AMUX_EN_VDDIO_H AMUX_EN_VDDIO_H_N AMUX_EN_VSWITCH_H
+ AMUX_EN_VSWITCH_H_N net74 ENABLE_VSWITCH_H VSSA VSWITCH
+ sky130_fd_io__gpiov2_amux_ctl_lshv2hv
Xpd_vdda_ls_q0 AMUX_EN_VDDIO_H AMUX_EN_VDDIO_H_N AMUX_EN_VDDA_H AMUX_EN_VDDA_H_N
+ ENABLE_VDDA_H_N ENABLE_VDDA_H VSSA VDDA sky130_fd_io__gpiov2_amux_ctl_lshv2hv
XI15 ANALOG_EN ana_en_i_n VSSD VCCD sky130_fd_io__gpiov2_amux_ctl_inv_1
XI16 ana_en_i_n ana_en_i VSSD VCCD sky130_fd_io__gpiov2_amux_ctl_inv_1
XI18 ENABLE_VSWITCH_H net74 VSSA VSWITCH sky130_fd_io__hvsbt_inv_x1
Xpd_vddio_ls_q0 ana_en_i ana_en_i_n AMUX_EN_VDDIO_H AMUX_EN_VDDIO_H_N HLD_I_H
+ HLD_I_H_N VSSD VDDIO_Q VCCD sky130_fd_io__gpiov2_amux_ctl_ls
.ENDS sky130_fd_io__gpiov2_amux_ls

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_ls_i2c_fix AMUX_EN_VDDA_H AMUX_EN_VDDA_H_N
+ AMUX_EN_VDDIO_H AMUX_EN_VSWITCH_H AMUX_EN_VSWITCH_H_N ANALOG_EN ENABLE_VDDA_H
+ ENABLE_VDDA_H_N ENABLE_VSWITCH_H HLD_I_H_N VCCD VDDA VDDIO_Q VSSA VSSD VSWITCH
*.PININFO AMUX_EN_VDDA_H:O AMUX_EN_VDDA_H_N:O AMUX_EN_VDDIO_H:O
*.PININFO AMUX_EN_VSWITCH_H:O AMUX_EN_VSWITCH_H_N:O ANALOG_EN:I
*.PININFO ENABLE_VDDA_H:I ENABLE_VDDA_H_N:O ENABLE_VSWITCH_H:I
*.PININFO HLD_I_H_N:I VCCD:I VDDA:I VDDIO_Q:I VSSA:I VSSD:I VSWITCH:I
Xpd_vddio_ls_q0 ana_en_i ana_en_i_n AMUX_EN_VDDIO_H net082 HLD_I_H_N VSSD
+ VDDIO_Q VCCD sky130_fd_io__gpiov2_amux_ctl_ls_i2c_fix
XI32 ENABLE_VDDA_H ENABLE_VDDA_H_N VSSA VDDA sky130_fd_io__gpiov2_amux_ls_inv_x1
Xpd_vswitch_ls_q0 AMUX_EN_VDDIO_H net028 AMUX_EN_VSWITCH_H AMUX_EN_VSWITCH_H_N
+ net83 ENABLE_VSWITCH_H VSSA VSWITCH sky130_fd_io__gpiov2_amux_ctl_lshv2hv
Xpd_vdda_ls_q0 AMUX_EN_VDDIO_H net028 AMUX_EN_VDDA_H AMUX_EN_VDDA_H_N
+ ENABLE_VDDA_H_N ENABLE_VDDA_H VSSA VDDA sky130_fd_io__gpiov2_amux_ctl_lshv2hv
XI15 ANALOG_EN ana_en_i_n VSSD VCCD sky130_fd_io__gpiov2_amux_ctl_inv_1
XI16 ana_en_i_n ana_en_i VSSD VCCD sky130_fd_io__gpiov2_amux_ctl_inv_1
XI18 ENABLE_VSWITCH_H net83 VSSA VSWITCH sky130_fd_io__hvsbt_inv_x1
XI36 AMUX_EN_VDDIO_H net028 VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
XI35 HLD_I_H_N net082 VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
.ENDS sky130_fd_io__gpiov2_amux_ls_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_ls_inv_x1 IN OUT VGND VPWR
*.PININFO IN:I OUT:O VGND:I VPWR:I
XI2 OUT IN VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.5 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amux_ls_inv_x1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_nand4 IN0 IN1 IN2 IN3 OUT VGND VPWR
*.PININFO IN0:I IN1:I IN2:I IN3:I OUT:O VGND:I VPWR:I
XI3 OUT IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI19 out_n OUT VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI20 OUT out_n VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN1 net50 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 net58 IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI15 net54 IN3 net58 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI14 net50 IN2 net54 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI18 out_n OUT VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI21 VGND out_n VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amux_nand4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_nand5 IN0 IN1 IN2 IN3 IN4 OUT VGND VPWR
*.PININFO IN0:I IN1:I IN2:I IN3:I IN4:I OUT:O VGND:I VPWR:I
XI3 OUT IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI20 OUT out_n VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI21 out_n OUT VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN1 net51 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI18 net63 IN4 net59 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 net59 IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI15 net55 IN3 net63 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI14 net51 IN2 net55 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI22 out_n OUT VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI23 VGND out_n VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amux_nand5

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amux_switch AMUXBUS_HV NG_AMX_VPMP_H NG_PAD_VPMP_H
+ NMID_VCCD PAD_HV_N0 PAD_HV_N1 PAD_HV_N2 PAD_HV_N3 PAD_HV_P0 PAD_HV_P1 PD_H_VDDA
+ PD_H_VDDIO PG_AMX_VDDA_H_N PG_PAD_VDDIOQ_H_N VDDA VDDIO VSSA VSSD
*.PININFO AMUXBUS_HV:B NG_AMX_VPMP_H:I NG_PAD_VPMP_H:I NMID_VCCD:I
*.PININFO PAD_HV_N0:B PAD_HV_N1:B PAD_HV_N2:B PAD_HV_N3:B PAD_HV_P0:B
*.PININFO PAD_HV_P1:B PD_H_VDDA:I PD_H_VDDIO:I PG_AMX_VDDA_H_N:I
*.PININFO PG_PAD_VDDIOQ_H_N:I VDDA:I VDDIO:I VSSA:I VSSD:I
xI72 VSSA VDDA sky130_fd_io__condiode
xI71 mid1 VDDA sky130_fd_io__condiode
xI70 mid VDDA sky130_fd_io__condiode
XI56 VSSA net79 sky130_fd_io__res75only_small
XI12 VSSA net77 sky130_fd_io__res75only_small
XI46 PAD_HV_N3 NG_PAD_VPMP_H mid1 mid1 sky130_fd_pr__nfet_g5v0d10v5 m=4 w=7.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI35 mid NG_PAD_VPMP_H PAD_HV_N1 mid sky130_fd_pr__nfet_g5v0d10v5 m=4 w=7.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI24 PAD_HV_N0 NG_PAD_VPMP_H mid mid sky130_fd_pr__nfet_g5v0d10v5 m=3 w=7.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI45 mid1 NG_PAD_VPMP_H PAD_HV_N2 mid1 sky130_fd_pr__nfet_g5v0d10v5 m=4 w=7.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI28 mid NG_AMX_VPMP_H AMUXBUS_HV mid sky130_fd_pr__nfet_g5v0d10v5 m=7 w=7.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI57 mid1 NMID_VCCD net79 VSSA sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI47 mid1 NG_AMX_VPMP_H AMUXBUS_HV mid1 sky130_fd_pr__nfet_g5v0d10v5 m=7 w=7.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI78<1> mid PD_H_VDDA VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI78<0> mid1 PD_H_VDDA VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI77<1> mid PD_H_VDDIO VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI77<0> mid1 PD_H_VDDIO VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 mid NMID_VCCD net77 VSSA sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI26 mid PG_AMX_VDDA_H_N AMUXBUS_HV VDDA sky130_fd_pr__pfet_g5v0d10v5 m=5 w=7.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI22 mid PG_PAD_VDDIOQ_H_N PAD_HV_P1 VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=3
+ w=7.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI36 mid PG_PAD_VDDIOQ_H_N PAD_HV_P0 VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=3
+ w=7.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
.ENDS sky130_fd_io__gpiov2_amux_switch

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amx_inv4 A Y VDA VSSA
*.PININFO A:I Y:O VDA:I VSSA:I
XI75 Y A VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=2 w=0.42 l=0.6 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI74 Y A VDA VDA sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amx_inv4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amx_pdcsd_inv A Y VDA VSSA
*.PININFO A:I Y:O VDA:I VSSA:I
XI414 Y A VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI519 Y VSSA VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI517 Y A VDA VDA sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=2.0 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI429 Y A VDA VDA sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.75 l=2.0 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amx_pdcsd_inv

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amx_pucsd_buf A Y VDA VSSA
*.PININFO A:I Y:O VDA:I VSSA:I
XI75 int A VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=4 w=0.42 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 Y int VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=3 w=0.42 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI74 int A VDA VDA sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI5 Y int VDA VDA sky130_fd_pr__pfet_g5v0d10v5 m=5 w=1.0 l=0.6 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amx_pucsd_buf

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_amx_pucsd_inv A Y VDA VSSA
*.PININFO A:I Y:O VDA:I VSSA:I
XI75 Y A VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 m=7 w=0.42 l=0.6 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI74 Y A VDA VDA sky130_fd_pr__pfet_g5v0d10v5 m=7 w=1.0 l=0.6 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_amx_pucsd_inv

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_ctl DM[2] DM[1] DM[0] DM_H[2] DM_H[1] DM_H[0]
+ DM_H_N[2] DM_H_N[1] DM_H_N[0] ENABLE_H ENABLE_INP_H HLD_H_N HLD_I_H HLD_I_H_N
+ HLD_I_OVR_H HLD_OVR IB_MODE_SEL IB_MODE_SEL_H IB_MODE_SEL_H_N INP_DIS
+ INP_DIS_H_N OD_I_H VCC_IO VGND VPWR VTRIP_SEL VTRIP_SEL_H VTRIP_SEL_H_N
*.PININFO DM[2]:I DM[1]:I DM[0]:I DM_H[2]:O DM_H[1]:O DM_H[0]:O
*.PININFO DM_H_N[2]:O DM_H_N[1]:O DM_H_N[0]:O ENABLE_H:I
*.PININFO ENABLE_INP_H:I HLD_H_N:I HLD_I_H:O HLD_I_H_N:O HLD_I_OVR_H:O
*.PININFO HLD_OVR:I IB_MODE_SEL:I IB_MODE_SEL_H:O IB_MODE_SEL_H_N:O
*.PININFO INP_DIS:I INP_DIS_H_N:O OD_I_H:O VCC_IO:I VGND:I VPWR:I
*.PININFO VTRIP_SEL:I VTRIP_SEL_H:O VTRIP_SEL_H_N:O
XI75 ENABLE_INP_H ENABLE_H startup_rst_h VGND VCC_IO sky130_fd_io__hvsbt_nor
Xhld_dis_blk_q0 ENABLE_H HLD_H_N HLD_I_H HLD_I_H_N HLD_I_OVR_H HLD_OVR OD_I_H
+ VCC_IO VGND VPWR sky130_fd_io__gpiov2_ctl_hld
Xls_bank_q0 DM[2] DM[1] DM[0] DM_H[2] DM_H[1] DM_H[0] DM_H_N[2] DM_H_N[1]
+ DM_H_N[0] HLD_I_H_N IB_MODE_SEL IB_MODE_SEL_H IB_MODE_SEL_H_N INP_DIS net80
+ INP_DIS_H_N OD_I_H startup_rst_h inp_startup_en_h VCC_IO VGND VPWR VTRIP_SEL
+ VTRIP_SEL_H VTRIP_SEL_H_N sky130_fd_io__gpiov2_ctl_lsbank
XI56 OD_I_H ENABLE_INP_H net92 VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI57 net92 inp_startup_en_h VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
.ENDS sky130_fd_io__gpiov2_ctl

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_ctl_hld ENABLE_H HLD_H_N HLD_I_H HLD_I_H_N
+ HLD_I_OVR_H HLD_OVR OD_I_H VCC_IO VGND VPWR
*.PININFO ENABLE_H:I HLD_H_N:I HLD_I_H:O HLD_I_H_N:O HLD_I_OVR_H:O
*.PININFO HLD_OVR:I OD_I_H:O VCC_IO:I VGND:I VPWR:I
Xhld_ovr_ls_q0 net65 HLD_OVR hld_ovr_h net37 od_h VGND VCC_IO VGND VPWR
+ sky130_fd_io__com_ctl_ls
XI30 OD_I_H hld_i_ovr_h_n HLD_I_OVR_H VGND VCC_IO sky130_fd_io__hvsbt_nor
XI26 net65 hld_ovr_h hld_i_ovr_h_n VGND VCC_IO sky130_fd_io__hvsbt_nor
Xhld_i_h_inv4_q0 net65 enable_vdda_h_n VGND VCC_IO sky130_fd_io__hvsbt_inv_x4
XI31 od_i_h_n OD_I_H VGND VCC_IO sky130_fd_io__hvsbt_inv_x4
Xhld_nand_q0 ENABLE_H HLD_H_N net64 VGND VCC_IO sky130_fd_io__hvsbt_nand2
Xod_h_inv_q0 ENABLE_H od_h VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
Xhld_i_h_inv1_q0 net64 net65 VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
XI32 od_h od_i_h_n VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
Xhld_i_h_inv8<1>_q0 enable_vdda_h_n hld_i_h_n_net<1> VGND VCC_IO
+ sky130_fd_io__hvsbt_inv_x8
Xhld_i_h_inv8<0>_q0 enable_vdda_h_n hld_i_h_n_net<0> VGND VCC_IO
+ sky130_fd_io__hvsbt_inv_x8
* Rshort<1> hld_i_h_n_net<1> HLD_I_H_N short
* Rshort<0> hld_i_h_n_net<0> HLD_I_H_N short
* Rshort_hld_i_h enable_vdda_h_n HLD_I_H short
Rshort<1> hld_i_h_n_net<1> HLD_I_H_N sky130_fd_pr__res_generic_m1 L=1 W=1
Rshort<0> hld_i_h_n_net<0> HLD_I_H_N sky130_fd_pr__res_generic_m1 L=1 W=1
Rshort_hld_i_h enable_vdda_h_n HLD_I_H sky130_fd_pr__res_generic_m1 L=1 W=1
.ENDS sky130_fd_io__gpiov2_ctl_hld

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_ctl_lsbank DM[2] DM[1] DM[0] DM_H[2] DM_H[1]
+ DM_H[0] DM_H_N[2] DM_H_N[1] DM_H_N[0] HLD_I_H_N IB_MODE_SEL IB_MODE_SEL_H
+ IB_MODE_SEL_H_N INP_DIS INP_DIS_H INP_DIS_H_N OD_I_H STARTUP_RST_H STARTUP_ST_H
+ VCC_IO VGND VPWR VTRIP_SEL VTRIP_SEL_H VTRIP_SEL_H_N
*.PININFO DM[2]:I DM[1]:I DM[0]:I DM_H[2]:O DM_H[1]:O DM_H[0]:O
*.PININFO DM_H_N[2]:O DM_H_N[1]:O DM_H_N[0]:O HLD_I_H_N:I
*.PININFO IB_MODE_SEL:I IB_MODE_SEL_H:O IB_MODE_SEL_H_N:O INP_DIS:I
*.PININFO INP_DIS_H:O INP_DIS_H_N:O OD_I_H:I STARTUP_RST_H:I
*.PININFO STARTUP_ST_H:I VCC_IO:I VGND:I VPWR:I VTRIP_SEL:I
*.PININFO VTRIP_SEL_H:O VTRIP_SEL_H_N:O
Xtrip_sel_st_q0 trip_sel_st_h OD_I_H VGND sky130_fd_io__tk_opti
Xtrip_sel_rst_q0 trip_sel_rst_h VGND OD_I_H sky130_fd_io__tk_opti
Xie_n_rst_q0 ie_n_rst_h STARTUP_RST_H STARTUP_ST_H sky130_fd_io__tk_opti
Xie_n_st_q0 ie_n_st_h STARTUP_ST_H STARTUP_RST_H sky130_fd_io__tk_opti
XI338<1> dm_rst_h<0> STARTUP_ST_H STARTUP_RST_H sky130_fd_io__tk_opti
XI803<1> dm_st_h<1> OD_I_H VGND sky130_fd_io__tk_opti
XI802<1> dm_st_h<2> OD_I_H VGND sky130_fd_io__tk_opti
XI804<1> dm_rst_h<2> VGND OD_I_H sky130_fd_io__tk_opti
XI805<1> dm_rst_h<1> VGND OD_I_H sky130_fd_io__tk_opti
* NOTE:  This has the selectable open and short on metal2 instead of metal1
XI598 ib_mode_sel_st_h OD_I_H VGND sky130_fd_io__tk_optiB
* NOTE:  This has the selectable short on metal2 instead of metal1
XI597 ib_mode_sel_rst_h VGND OD_I_H sky130_fd_io__tk_optiA
XI337<1> dm_st_h<0> STARTUP_RST_H STARTUP_ST_H sky130_fd_io__tk_opti
Xdm_ls<0>_q0 HLD_I_H_N DM[0] DM_H[0] DM_H_N[0] dm_rst_h<0> dm_st_h<0> VCC_IO
+ VGND VPWR sky130_fd_io__com_ctl_ls
Xinp_dis_ls_q0 HLD_I_H_N INP_DIS INP_DIS_H INP_DIS_H_N ie_n_rst_h ie_n_st_h
+ VCC_IO VGND VPWR sky130_fd_io__com_ctl_ls
Xtrip_sel_ls_q0 HLD_I_H_N VTRIP_SEL VTRIP_SEL_H VTRIP_SEL_H_N trip_sel_rst_h
+ trip_sel_st_h VCC_IO VGND VPWR sky130_fd_io__com_ctl_ls
Xdm_ls<2>_q0 HLD_I_H_N DM[2] DM_H[2] DM_H_N[2] dm_rst_h<2> dm_st_h<2> VCC_IO
+ VGND VPWR sky130_fd_io__com_ctl_ls
Xdm_ls<1>_q0 HLD_I_H_N DM[1] DM_H[1] DM_H_N[1] dm_rst_h<1> dm_st_h<1> VCC_IO
+ VGND VPWR sky130_fd_io__com_ctl_ls
XI595 HLD_I_H_N IB_MODE_SEL IB_MODE_SEL_H IB_MODE_SEL_H_N ib_mode_sel_rst_h
+ ib_mode_sel_st_h VCC_IO VGND VPWR sky130_fd_io__com_ctl_ls
.ENDS sky130_fd_io__gpiov2_ctl_lsbank

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_ibuf_se ENABLE_VDDIO_LV IBUFMUX_OUT IBUFMUX_OUT_H
+ IN_H IN_VT MODE_NORMAL_N MODE_VCCHIB_N VCCHIB VDDIO_Q VSSD VTRIP_SEL_H
+ VTRIP_SEL_H_N
*.PININFO ENABLE_VDDIO_LV:I IBUFMUX_OUT:O IBUFMUX_OUT_H:O IN_H:I
*.PININFO IN_VT:I MODE_NORMAL_N:I MODE_VCCHIB_N:I VCCHIB:I VDDIO_Q:I
*.PININFO VSSD:I VTRIP_SEL_H:I VTRIP_SEL_H_N:I
XI148 ENABLE_VDDIO_LV mode_vcchib mode_vcchib_lv_n VSSD VCCHIB
+ sky130_fd_io__hvsbt_nand2
XI149 ENABLE_VDDIO_LV mode_normal mode_normal_lv_n VSSD VCCHIB
+ sky130_fd_io__hvsbt_nand2
XI112 mode_normal_lv_n mode_normal_lv VSSD VSSD VCCHIB VCCHIB
+ sky130_fd_io__gpiov2_inbuf_lvinv_x1
XI111 mode_vcchib_lv_n mode_vcchib_lv VSSD VSSD VCCHIB VCCHIB
+ sky130_fd_io__gpiov2_inbuf_lvinv_x1
Xlvls_q0 out_vcchib out_vddio mode_normal_lv mode_normal_lv_n mode_vcchib_lv
+ mode_vcchib_lv_n IBUFMUX_OUT net57 VCCHIB VSSD sky130_fd_io__gpiov2_ipath_lvls
Xhvls_q0 out_vcchib out_vddio out_n_vcchib mode_normal MODE_NORMAL_N mode_vcchib
+ MODE_VCCHIB_N IBUFMUX_OUT_H net68 VDDIO_Q VSSD sky130_fd_io__gpiov2_ipath_hvls
XI88 IN_H mode_vcchib_lv_n out_vcchib out_n_vcchib VCCHIB VSSD
+ sky130_fd_io__gpiov2_vcchib_in_buf
Xbuf_q0 IN_H IN_VT MODE_NORMAL_N out_vddio out_n_vddio VDDIO_Q VSSD VTRIP_SEL_H
+ VTRIP_SEL_H_N sky130_fd_io__gpiov2_in_buf
XI491 MODE_NORMAL_N mode_normal VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
XI105 MODE_VCCHIB_N mode_vcchib VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
.ENDS sky130_fd_io__gpiov2_ibuf_se

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_ictl_logic DM_H_N[2] DM_H_N[1] DM_H_N[0]
+ IB_MODE_SEL_H IB_MODE_SEL_H_N INP_DIS_H_N INP_DIS_I_H INP_DIS_I_H_N
+ MODE_NORMAL_N MODE_VCCHIB_N TRIPSEL_I_H TRIPSEL_I_H_N VDDIO_Q VSSD VTRIP_SEL_H_N
*.PININFO DM_H_N[2]:I DM_H_N[1]:I DM_H_N[0]:I IB_MODE_SEL_H:I
*.PININFO IB_MODE_SEL_H_N:I INP_DIS_H_N:I INP_DIS_I_H:O
*.PININFO INP_DIS_I_H_N:O MODE_NORMAL_N:O MODE_VCCHIB_N:O
*.PININFO TRIPSEL_I_H:O TRIPSEL_I_H_N:O VDDIO_Q:I VSSD:I
*.PININFO VTRIP_SEL_H_N:I
XI71 VTRIP_SEL_H_N MODE_NORMAL_N TRIPSEL_I_H VSSD VDDIO_Q
+ sky130_fd_io__hvsbt_nor
XI80 dm_buf_dis_n INP_DIS_H_N INP_DIS_I_H VSSD VDDIO_Q sky130_fd_io__hvsbt_nand2
XI79 DM_H_N[2] and_dm01 dm_buf_dis_n VSSD VDDIO_Q sky130_fd_io__hvsbt_nand2
XI78 DM_H_N[1] DM_H_N[0] nand_dm01 VSSD VDDIO_Q sky130_fd_io__hvsbt_nand2
XI36 INP_DIS_I_H_N IB_MODE_SEL_H MODE_VCCHIB_N VSSD VDDIO_Q
+ sky130_fd_io__hvsbt_nand2
XI35 INP_DIS_I_H_N IB_MODE_SEL_H_N MODE_NORMAL_N VSSD VDDIO_Q
+ sky130_fd_io__hvsbt_nand2
XI111 INP_DIS_I_H INP_DIS_I_H_N VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
XI75 nand_dm01 and_dm01 VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
XI74 TRIPSEL_I_H TRIPSEL_I_H_N VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
.ENDS sky130_fd_io__gpiov2_ictl_logic

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_in_buf IN_H IN_VT MODE_NORMAL_N OUT OUT_N VDDIO_Q
+ VSSD VTRIP_SEL_H VTRIP_SEL_H_N
*.PININFO IN_H:I IN_VT:I MODE_NORMAL_N:I OUT:O OUT_N:O VDDIO_Q:I
*.PININFO VSSD:I VTRIP_SEL_H:I VTRIP_SEL_H_N:I
XI43 mode_normal_cmos_h mode_normal_cmos_h_n VSSD VDDIO_Q
+ sky130_fd_io__hvsbt_inv_x1
XI488 VTRIP_SEL_H MODE_NORMAL_N mode_normal_cmos_h VSSD VDDIO_Q
+ sky130_fd_io__hvsbt_nor
XI583 IN_VT VTRIP_SEL_H_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI644 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI646 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI593 net91 MODE_NORMAL_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI592 net103 in_b fbk VSSD sky130_fd_pr__nfet_g5v0d10v5 m=4 w=1.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI591 fbk IN_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=6 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI590 fbk2 in_b fbk VSSD sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI589 net91 in_b VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI588 fbk IN_VT VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI587 in_b IN_H fbk VSSD sky130_fd_pr__nfet_g5v0d10v5 m=5 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI586 OUT_N net91 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI642 OUT OUT_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI629 in_b IN_H net158 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.8
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI636 net158 mode_normal_cmos_h_n VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5
+ m=2 w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI632 net122 MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=2
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI647 VDDIO_Q VDDIO_Q VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0
+ l=0.8 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI600 net103 MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=2
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI598 net91 in_b net138 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI597 fbk2 mode_normal_cmos_h_n VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=2
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI596 OUT_N net91 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI595 net138 MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI631 in_b IN_H net122 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.8
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI643 OUT OUT_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_in_buf

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_inbuf_lvinv_x1 IN OUT VGND VNB VPB VPWR
*.PININFO IN:I OUT:O VGND:I VNB:I VPB:I VPWR:I
XI2 OUT IN VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=1.0 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=3.0 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_inbuf_lvinv_x1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_ipath DM_H_N[2] DM_H_N[1] DM_H_N[0] ENABLE_VDDIO_LV
+ IB_MODE_SEL_H IB_MODE_SEL_H_N INP_DIS_H_N OUT OUT_H PAD VCCHIB VDDIO_Q VSSD
+ VTRIP_SEL_H_N
*.PININFO DM_H_N[2]:I DM_H_N[1]:I DM_H_N[0]:I ENABLE_VDDIO_LV:I
*.PININFO IB_MODE_SEL_H:I IB_MODE_SEL_H_N:I INP_DIS_H_N:I OUT:O
*.PININFO OUT_H:O PAD:B VCCHIB:I VDDIO_Q:I VSSD:I VTRIP_SEL_H_N:I
XI106 ENABLE_VDDIO_LV OUT OUT_H in_h in_vt mode_normal_n mode_vcchib_n VCCHIB
+ VDDIO_Q VSSD tripsel_i_h tripsel_i_h_n sky130_fd_io__gpiov2_ibuf_se
XI107 DM_H_N[2] DM_H_N[1] DM_H_N[0] IB_MODE_SEL_H IB_MODE_SEL_H_N INP_DIS_H_N
+ en_h_n en_h mode_normal_n mode_vcchib_n tripsel_i_h tripsel_i_h_n VDDIO_Q VSSD
+ VTRIP_SEL_H_N sky130_fd_io__gpiov2_ictl_logic
XI120 PAD in_h in_vt VDDIO_Q VSSD tripsel_i_h
+ sky130_fd_io__gpio_ovtv2_buf_localesd
.ENDS sky130_fd_io__gpiov2_ipath

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_ipath_hvls IN_VCCHIB IN_VDDIO INB_VCCHIB
+ MODE_NORMAL MODE_NORMAL_N MODE_VCCHIB MODE_VCCHIB_N OUT OUT_B VDDIO_Q VSSD
*.PININFO IN_VCCHIB:I IN_VDDIO:I INB_VCCHIB:I MODE_NORMAL:I
*.PININFO MODE_NORMAL_N:I MODE_VCCHIB:I MODE_VCCHIB_N:I OUT:O OUT_B:O
*.PININFO VDDIO_Q:I VSSD:I
XI325 fbk fbk_b VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI324 fbk_b fbk VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI323 net63 MODE_NORMAL VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI322 OUT_B IN_VDDIO net75 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI321 net75 MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI320 OUT OUT_B VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=5 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI319 OUT_B MODE_VCCHIB net63 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI318 net55 MODE_VCCHIB_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI317 OUT_B net84 net55 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI336 net84 fbk_b VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI335 OUT_B net84 net88 VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI334 fbk INB_VCCHIB net116 VSSD sky130_fd_pr__nfet_g5v0d10v5 m=3 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI333 net116 MODE_VCCHIB VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI332 net112 MODE_NORMAL VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI331 OUT OUT_B VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=3 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI330 OUT_B IN_VDDIO net112 VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI329 fbk_b IN_VCCHIB net92 VSSD sky130_fd_pr__nfet_g5v0d10v5 m=3 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI328 fbk MODE_VCCHIB_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI327 net92 MODE_VCCHIB VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI326 net88 MODE_VCCHIB VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI337 net84 fbk_b VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_ipath_hvls

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_ipath_lvls IN_VCCHIB IN_VDDIO MODE_NORMAL_LV
+ MODE_NORMAL_LV_N MODE_VCCHIB_LV MODE_VCCHIB_LV_N OUT OUT_B VCCHIB VSSD
*.PININFO IN_VCCHIB:I IN_VDDIO:I MODE_NORMAL_LV:I MODE_NORMAL_LV_N:I
*.PININFO MODE_VCCHIB_LV:I MODE_VCCHIB_LV_N:I OUT:O OUT_B:O VCCHIB:I
*.PININFO VSSD:I
XI345 fbk_n IN_VDDIO VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI344 net70 MODE_VCCHIB_LV VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 m=1 w=3.0
+ l=0.25 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI343 OUT_B fbk net78 VCCHIB sky130_fd_pr__pfet_01v8 m=2 w=3.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI342 net78 MODE_NORMAL_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 m=2 w=3.0
+ l=0.25 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI341 OUT_B MODE_NORMAL_LV net70 VCCHIB sky130_fd_pr__pfet_01v8 m=1 w=3.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI340 net50 MODE_VCCHIB_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 m=2 w=3.0
+ l=0.25 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI339 fbk_n MODE_NORMAL_LV VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 m=1 w=5.0
+ l=0.25 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI338 fbk fbk_n VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 m=1 w=5.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI337 OUT OUT_B VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 m=4 w=3.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI336 OUT_B IN_VCCHIB net50 VCCHIB sky130_fd_pr__pfet_01v8 m=2 w=3.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI351 net111 MODE_NORMAL_LV VSSD VSSD sky130_fd_pr__nfet_01v8 m=2 w=3.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI350 OUT_B fbk net111 VSSD sky130_fd_pr__nfet_01v8 m=2 w=3.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI349 OUT OUT_B VSSD VSSD sky130_fd_pr__nfet_01v8 m=2 w=3.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI348 fbk fbk_n VSSD VSSD sky130_fd_pr__nfet_01v8 m=1 w=3.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI347 net95 MODE_VCCHIB_LV VSSD VSSD sky130_fd_pr__nfet_01v8 m=2 w=3.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI346 OUT_B IN_VCCHIB net95 VSSD sky130_fd_pr__nfet_01v8 m=2 w=3.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI353 fbk_n IN_VDDIO net115 VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI352 net115 MODE_NORMAL_LV VSSD VSSD sky130_fd_pr__nfet_01v8 m=1 w=3.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_ipath_lvls

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_obpredrvr DRVHI_H DRVLO_H_N I2C_MODE_H_N PD_H[4]
+ PD_H[3] PD_H[2] PD_H[1] PD_H[0] PDEN_H_N[1] PDEN_H_N[0] PU_H_N[3] PU_H_N[2]
+ PU_H_N[1] PU_H_N[0] PUEN_H[1] PUEN_H[0] SLOW_H SLOW_H_N TIE_HI_ESD VCC_IO VGND
+ VGND_IO
*.PININFO DRVHI_H:I DRVLO_H_N:I I2C_MODE_H_N:I PD_H[4]:O PD_H[3]:O
*.PININFO PD_H[2]:O PD_H[1]:O PD_H[0]:O PDEN_H_N[1]:I PDEN_H_N[0]:I
*.PININFO PU_H_N[3]:O PU_H_N[2]:O PU_H_N[1]:O PU_H_N[0]:O PUEN_H[1]:I
*.PININFO PUEN_H[0]:I SLOW_H:I SLOW_H_N:I TIE_HI_ESD:I VCC_IO:I VGND:I
*.PININFO VGND_IO:I
Xpu_strong_q0 DRVHI_H PU_H_N[3] PU_H_N[2] PUEN_H[1] SLOW_H_N VCC_IO VGND_IO
+ sky130_fd_io__gpiov2_pupredrvr_strong
Xpd_strong_q0 DRVLO_H_N I2C_MODE_H_N PD_H[4] PD_H[3] PD_H[2] PDEN_H_N[1] SLOW_H
+ TIE_HI_ESD VCC_IO VGND VGND_IO sky130_fd_io__gpiov2_pdpredrvr_strong
Xpu_weak_q0 DRVHI_H PU_H_N[0] PUEN_H[0] VCC_IO VGND_IO
+ sky130_fd_io__com_pupredrvr_weak
Xpd_weak_q0 DRVLO_H_N PD_H[0] PDEN_H_N[0] VCC_IO VGND_IO
+ sky130_fd_io__com_pdpredrvr_weak
Xpu_strong_slow_q0 DRVHI_H PU_H_N[1] PUEN_H[1] VCC_IO VGND_IO
+ sky130_fd_io__com_pupredrvr_strong_slow
Xpd_strong_slow_q0 DRVLO_H_N PD_H[1] PDEN_H_N[1] VCC_IO VGND_IO
+ sky130_fd_io__com_pdpredrvr_strong_slow
xI15 VGND_IO VCC_IO sky130_fd_io__condiode
.ENDS sky130_fd_io__gpiov2_obpredrvr

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_octl DM_H[2] DM_H[1] DM_H[0] DM_H_N[2] DM_H_N[1]
+ DM_H_N[0] HLD_I_H_N OD_H PDEN_H_N[2] PDEN_H_N[1] PDEN_H_N[0] PUEN_0_H
+ PUEN_2OR1_H PUEN_H[1] PUEN_H[0] SLOW SLOW_H SLOW_H_N VCC_IO VGND VPWR
+ VREG_EN_H_N
*.PININFO DM_H[2]:I DM_H[1]:I DM_H[0]:I DM_H_N[2]:I DM_H_N[1]:I
*.PININFO DM_H_N[0]:I HLD_I_H_N:I OD_H:I PDEN_H_N[2]:O PDEN_H_N[1]:O
*.PININFO PDEN_H_N[0]:O PUEN_0_H:O PUEN_2OR1_H:O PUEN_H[1]:O
*.PININFO PUEN_H[0]:O SLOW:I SLOW_H:O SLOW_H_N:O VCC_IO:I VGND:I
*.PININFO VPWR:I VREG_EN_H_N:I
XI211 n<8> DM_H_N[1] PUEN_0_H VGND VCC_IO sky130_fd_io__hvsbt_nor
XI201 DM_H_N[2] DM_H_N[1] n<9> VGND VCC_IO sky130_fd_io__hvsbt_nor
XI381 DM_H[1] DM_H[0] net70 VGND VCC_IO sky130_fd_io__hvsbt_nor
XI210 DM_H[2] DM_H[0] n<8> VGND VCC_IO sky130_fd_io__hvsbt_xor
XI200 DM_H[2] DM_H[1] n<10> VGND VCC_IO sky130_fd_io__hvsbt_xor
XI185 DM_H_N[0] n<4> net130 VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI186 DM_H_N[2] DM_H_N[1] n<4> VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI187 DM_H[1] DM_H[0] n<3> VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI208 PUEN_2OR1_H VREG_EN_H_N n<5> VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI203 n<10> DM_H[0] n<1> VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI204 n<9> DM_H_N[0] n<0> VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI205 n<1> n<0> PUEN_2OR1_H VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI382 DM_H[2] net70 PDEN_H_N[2] VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI254 puen_h1_n PUEN_H[1] VGND VCC_IO sky130_fd_io__hvsbt_inv_x2
XI256 puen_h0_n PUEN_H[0] VGND VCC_IO sky130_fd_io__hvsbt_inv_x2
XI249 pden_h0 PDEN_H_N[0] VGND VCC_IO sky130_fd_io__hvsbt_inv_x2
XI247 pden_h1 PDEN_H_N[1] VGND VCC_IO sky130_fd_io__hvsbt_inv_x2
XI377 PUEN_0_H puen_h0_n VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
XI209 n<5> n<2> VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
XI376 n<2> puen_h1_n VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
XI374 net130 pden_h1 VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
XI375 n<3> pden_h0 VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
Xls_slow_q0 HLD_I_H_N SLOW SLOW_H SLOW_H_N OD_H VGND VCC_IO VGND VPWR
+ sky130_fd_io__com_ctl_ls
.ENDS sky130_fd_io__gpiov2_octl

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_octl_dat DM_H[2] DM_H[1] DM_H[0] DM_H_N[2]
+ DM_H_N[1] DM_H_N[0] DRVHI_H HLD_I_H_N HLD_I_OVR_H OD_H OE_N OUT PD_H[4] PD_H[3]
+ PD_H[2] PD_H[1] PD_H[0] PU_H_N[3] PU_H_N[2] PU_H_N[1] PU_H_N[0] SLOW SLOW_H_N
+ TIE_HI_ESD VCC_IO VGND VGND_IO VPWR VPWR_KA
*.PININFO DM_H[2]:I DM_H[1]:I DM_H[0]:I DM_H_N[2]:I DM_H_N[1]:I
*.PININFO DM_H_N[0]:I DRVHI_H:O HLD_I_H_N:I HLD_I_OVR_H:I OD_H:I
*.PININFO OE_N:I OUT:I PD_H[4]:O PD_H[3]:O PD_H[2]:O PD_H[1]:O
*.PININFO PD_H[0]:O PU_H_N[3]:O PU_H_N[2]:O PU_H_N[1]:O PU_H_N[0]:O
*.PININFO SLOW:I SLOW_H_N:O TIE_HI_ESD:I VCC_IO:I VGND:I VGND_IO:I
*.PININFO VPWR:I VPWR_KA:I
Xdatoe_q0 DRVHI_H drvlo_h_n HLD_I_H_N HLD_I_OVR_H OD_H oe_h OE_N OUT VCC_IO VGND
+ VPWR_KA sky130_fd_io__gpiov2_opath_datoe
Xctl_q0 DM_H[2] DM_H[1] DM_H[0] DM_H_N[2] DM_H_N[1] DM_H_N[0] HLD_I_H_N OD_H
+ pden_h_n<2> pden_h_n<1> pden_h_n<0> puen_0_h puen_2or1_h puen_h<1> puen_h<0>
+ SLOW slow_h SLOW_H_N VCC_IO VGND VPWR VCC_IO sky130_fd_io__gpiov2_octl
Xpredrvr_q0 DRVHI_H drvlo_h_n pden_h_n<2> PD_H[4] PD_H[3] PD_H[2] PD_H[1]
+ PD_H[0] pden_h_n<1> pden_h_n<0> PU_H_N[3] PU_H_N[2] PU_H_N[1] PU_H_N[0]
+ puen_h<1> puen_h<0> slow_h SLOW_H_N TIE_HI_ESD VCC_IO VGND VGND_IO
+ sky130_fd_io__gpiov2_obpredrvr
.ENDS sky130_fd_io__gpiov2_octl_dat

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_octl_mux A_H B_H SEL_H SEL_H_N VCCIO VSSIO Y_H
*.PININFO A_H:I B_H:I SEL_H:I SEL_H_N:I VCCIO:I VSSIO:I Y_H:O
XI2 Y_H SEL_H B_H VCCIO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI3 Y_H SEL_H_N A_H VCCIO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 B_H SEL_H_N Y_H VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI4 A_H SEL_H Y_H VSSIO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_octl_mux

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_odrvr FORCE_HI_H_N PAD PD_H[3] PD_H[2] PD_H[1]
+ PD_H[0] PD_H_I2C PU_H_N[3] PU_H_N[2] PU_H_N[1] PU_H_N[0] TIE_HI_ESD TIE_LO_ESD
+ VCC_IO VGND VGND_IO
*.PININFO FORCE_HI_H_N:I PAD:O PD_H[3]:I PD_H[2]:I PD_H[1]:I PD_H[0]:I
*.PININFO PD_H_I2C:I PU_H_N[3]:I PU_H_N[2]:I PU_H_N[1]:I PU_H_N[0]:I
*.PININFO TIE_HI_ESD:O TIE_LO_ESD:O VCC_IO:I VGND:I VGND_IO:I
Xodrvr_q0 FORCE_HI_H_N PAD PD_H[3] PD_H[2] PD_H[1] PD_H[0] PD_H_I2C PU_H_N[3]
+ PU_H_N[2] PU_H_N[1] PU_H_N[0] TIE_HI_ESD TIE_LO_ESD VCC_IO VGND VGND_IO
+ sky130_fd_io__gpiov2_odrvr_sub
Xbondpad_q0 PAD VGND_IO sky130_fd_io__com_pad
.ENDS sky130_fd_io__gpiov2_odrvr

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_odrvr_sub FORCE_HI_H_N PAD PD_H[3] PD_H[2] PD_H[1]
+ PD_H[0] PD_H_I2C PU_H_N[3] PU_H_N[2] PU_H_N[1] PU_H_N[0] TIE_HI_ESD TIE_LO_ESD
+ VCC_IO VGND VGND_IO
*.PININFO FORCE_HI_H_N:I PAD:O PD_H[3]:I PD_H[2]:I PD_H[1]:I PD_H[0]:I
*.PININFO PD_H_I2C:I PU_H_N[3]:I PU_H_N[2]:I PU_H_N[1]:I PU_H_N[0]:I
*.PININFO TIE_HI_ESD:B TIE_LO_ESD:B VCC_IO:I VGND:I VGND_IO:I
Xpddrvr_strong_q0 PAD PD_H[3] PD_H[2] PD_H_I2C TIE_LO_ESD VCC_IO VGND_IO
+ sky130_fd_io__gpiov2_pddrvr_strong
Xpudrvr_strong_q0 PAD PU_H_N[3] PU_H_N[2] TIE_HI_ESD VCC_IO VGND
+ sky130_fd_io__gpio_pudrvr_strong
Xpudrvr_weak_q0 weak_pad PU_H_N[0] VCC_IO VGND VCC_IO
+ sky130_fd_io__com_pudrvr_weak
Xpddrvr_weak_q0 weak_pad PD_H[0] VCC_IO VGND_IO sky130_fd_io__gpio_pddrvr_weak
Xstrong_slow_pddrvr_q0 strong_slow_pad PD_H[1] VCC_IO VGND_IO
+ sky130_fd_io__gpio_pddrvr_strong_slow
Xstrong_slow_pudrvr_q0 strong_slow_pad PU_H_N[1] VCC_IO VGND VCC_IO
+ sky130_fd_io__com_pudrvr_strong_slow
Xres_q0 strong_slow_pad pad_r250 VGND_IO sky130_fd_io__com_res_strong_slow
Xres_weak_q0 weak_pad pad_r250 VGND_IO sky130_fd_io__com_res_weak
Xresd_q0 PAD pad_r250 sky130_fd_io__res250only_small
xI60 VGND_IO VCC_IO sky130_fd_io__condiode
xI59 VGND_IO VCC_IO sky130_fd_io__condiode
xI58 VGND_IO VCC_IO sky130_fd_io__condiode
xI72 VGND_IO VCC_IO sky130_fd_io__condiode
.ENDS sky130_fd_io__gpiov2_odrvr_sub

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_opath DM_H[2] DM_H[1] DM_H[0] DM_H_N[2] DM_H_N[1]
+ DM_H_N[0] HLD_I_H_N HLD_I_OVR_H OD_H OE_N OUT PAD SLOW TIE_HI_ESD TIE_LO_ESD
+ VCC_IO VGND VGND_IO VPWR VPWR_KA
*.PININFO DM_H[2]:I DM_H[1]:I DM_H[0]:I DM_H_N[2]:I DM_H_N[1]:I
*.PININFO DM_H_N[0]:I HLD_I_H_N:I HLD_I_OVR_H:I OD_H:I OE_N:I OUT:I
*.PININFO PAD:O SLOW:I TIE_HI_ESD:O TIE_LO_ESD:O VCC_IO:I VGND:I
*.PININFO VGND_IO:I VPWR:I VPWR_KA:I
Xodrvr_q0 net70 PAD pd_h<3> pd_h<2> pd_h<1> pd_h<0> pd_h<4> pu_h_n<3> pu_h_n<2>
+ pu_h_n<1> pu_h_n<0> TIE_HI_ESD TIE_LO_ESD VCC_IO VGND VGND_IO
+ sky130_fd_io__gpiov2_odrvr
Xopath_q0 DM_H[2] DM_H[1] DM_H[0] DM_H_N[2] DM_H_N[1] DM_H_N[0] drvhi_h
+ HLD_I_H_N HLD_I_OVR_H OD_H OE_N OUT pd_h<4> pd_h<3> pd_h<2> pd_h<1> pd_h<0>
+ pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> SLOW slow_h_n TIE_HI_ESD VCC_IO VGND
+ VGND_IO VPWR VPWR_KA sky130_fd_io__gpiov2_octl_dat
.ENDS sky130_fd_io__gpiov2_opath

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_opath_datoe DRVHI_H DRVLO_H_N HLD_H_N HLD_I_OVR_H
+ OD_H OE_H OE_N OUT VCC_IO VGND VPWR_KA
*.PININFO DRVHI_H:O DRVLO_H_N:O HLD_H_N:I HLD_I_OVR_H:I OD_H:I OE_H:O
*.PININFO OE_N:I OUT:I VCC_IO:I VGND:I VPWR_KA:I
Xdat_ls_q0 HLD_I_OVR_H OUT pd_dis_h pu_dis_h VGND OD_H VCC_IO VGND VPWR_KA
+ sky130_fd_io__gpio_dat_ls
Xoe_ls_q0 HLD_I_OVR_H OE_N oe_h_n OE_H VGND OD_H VCC_IO VGND VPWR_KA
+ sky130_fd_io__gpio_dat_ls
Xcclat_q0 DRVHI_H DRVLO_H_N oe_h_n pd_dis_h pu_dis_h VCC_IO VGND
+ sky130_fd_io__com_cclat
.ENDS sky130_fd_io__gpiov2_opath_datoe

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_pddrvr_strong PAD PD_H[3] PD_H[2] PD_H_I2C
+ TIE_LO_ESD VCC_IO VGND_IO
*.PININFO PAD:O PD_H[3]:I PD_H[2]:I PD_H_I2C:I TIE_LO_ESD:O VCC_IO:I
*.PININFO VGND_IO:I
XI97 PD_H[3] net80 sky130_fd_io__tk_em2s
XI108 PD_H[3] net78 sky130_fd_io__tk_em2s
XI109 TIE_LO_ESD net76 sky130_fd_io__tk_em2s
XI102 PD_H[3] net72 sky130_fd_io__tk_em2s
XI104 PD_H[3] net68 sky130_fd_io__tk_em2s
XI96 PD_H[3] net66 sky130_fd_io__tk_em2s
XI113 PD_H[2] net46 sky130_fd_io__tk_em2s
XI99 TIE_LO_ESD net80 sky130_fd_io__tk_em2o
XI98 PD_H[2] net80 sky130_fd_io__tk_em2o
XI106 PD_H[2] net78 sky130_fd_io__tk_em2o
XI107 TIE_LO_ESD net78 sky130_fd_io__tk_em2o
XI110 PD_H[3] net76 sky130_fd_io__tk_em2o
XI111 PD_H[2] net76 sky130_fd_io__tk_em2o
XI100 TIE_LO_ESD net72 sky130_fd_io__tk_em2o
XI101 PD_H[2] net72 sky130_fd_io__tk_em2o
XI103 TIE_LO_ESD net68 sky130_fd_io__tk_em2o
XI105 PD_H[2] net68 sky130_fd_io__tk_em2o
XI95 PD_H[2] net66 sky130_fd_io__tk_em2o
XI94 TIE_LO_ESD net66 sky130_fd_io__tk_em2o
XI88 PD_H[3] net46 sky130_fd_io__tk_em2o
XI87 TIE_LO_ESD net46 sky130_fd_io__tk_em2o
XI49 VGND_IO TIE_LO_ESD sky130_fd_io__tk_tie_r_out_esd
Xn24<2>_q0 PAD net80 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn24<1>_q0 PAD net80 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn24<0>_q0 PAD net80 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn23<2>_q0 PAD net66 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn23<1>_q0 PAD net66 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn23<0>_q0 PAD net66 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn22<2>_q0 PAD PD_H[3] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn22<1>_q0 PAD PD_H[3] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn22<0>_q0 PAD PD_H[3] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn21<2>_q0 PAD PD_H[3] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn21<1>_q0 PAD PD_H[3] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn21<0>_q0 PAD PD_H[3] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn12_q0 PAD PD_H_I2C VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn32<2>_q0 PAD net68 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn32<1>_q0 PAD net68 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn32<0>_q0 PAD net68 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn33<2>_q0 PAD net78 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn33<1>_q0 PAD net78 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn33<0>_q0 PAD net78 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn34<3>_q0 PAD net76 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn34<2>_q0 PAD net76 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn34<1>_q0 PAD net76 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn34<0>_q0 PAD net76 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn11<2>_q0 PAD PD_H[2] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn11<1>_q0 PAD PD_H[2] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn11<0>_q0 PAD PD_H[2] VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn13_q0 PAD net46 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
Xn31_q0 PAD net72 VGND_IO sky130_fd_io__com_pddrvr_unit_2_5
xI72 VGND_IO VCC_IO sky130_fd_io__condiode
.ENDS sky130_fd_io__gpiov2_pddrvr_strong

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_pdpredrvr_strong DRVLO_H_N I2C_MODE_H_N PD_H[4]
+ PD_H[3] PD_H[2] PDEN_H_N SLOW_H TIE_HI_ESD VCC_IO VGND VGND_IO
*.PININFO DRVLO_H_N:I I2C_MODE_H_N:I PD_H[4]:O PD_H[3]:O PD_H[2]:O
*.PININFO PDEN_H_N:I SLOW_H:I TIE_HI_ESD:I VCC_IO:I VGND:I VGND_IO:I
XI160 I2C_MODE_H_N SLOW_H net75 VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI98 i2c_mode_h SLOW_H int_slow1 VGND VCC_IO sky130_fd_io__hvsbt_nand2
XI161 net75 net142 VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
XI97 int_slow1 mod_slow_h VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
XI93 I2C_MODE_H_N i2c_mode_h VGND VCC_IO sky130_fd_io__hvsbt_inv_x1
Xmux_q0 mod_drvlo_h_n_i2c DRVLO_H_N i2c_mode_h I2C_MODE_H_N VCC_IO VGND_IO
+ mod_drvlo_h_n sky130_fd_io__gpiov2_octl_mux
Xnr3_q0 DRVLO_H_N pbias_out pbias_out mod_slow_h PD_H[2] PD_H[4] PDEN_H_N VCC_IO
+ VGND_IO sky130_fd_io__gpiov2_pdpredrvr_strong_nr2
Xnr2_q0 mod_drvlo_h_n en_fast2_n<1> en_fast2_n<0> mod_slow_h PD_H[3] PDEN_H_N
+ VCC_IO VGND_IO sky130_fd_io__gpiov2_pdpredrvr_strong_nr3
XI77 en_fast2_n<1> pbias_out en_fast_h_n sky130_fd_io__tk_opto
XI76 net118 pbias_out en_fast_h_n sky130_fd_io__tk_opto
XI79 en_fast2_n<0> en_fast2_n<1> VCC_IO sky130_fd_io__tk_opti
Xinv_q0 en_fast_h en_fast_h_n VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
Xbias_q0 DRVLO_H_N en_fast_h en_fast_h_n pbias_out PD_H[4] PDEN_H_N VCC_IO
+ VGND_IO sky130_fd_io__com_pdpredrvr_pbias
Xnor_q0 net142 PDEN_H_N en_fast_h VGND_IO VCC_IO sky130_fd_io__com_nor2_dnw
XI87 mod_drvlo_h_n_i2c PD_H[4] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=3.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI88 mod_drvlo_h_n_i2c PD_H[4] VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_pdpredrvr_strong

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_pdpredrvr_strong_nr2 DRVLO_H_N EN_FAST_N[1]
+ EN_FAST_N[0] I2C_MODE_H PD_H PD_I2C_H PDEN_H_N VCC_IO VGND_IO
*.PININFO DRVLO_H_N:I EN_FAST_N[1]:I EN_FAST_N[0]:I I2C_MODE_H:I
*.PININFO PD_H:O PD_I2C_H:O PDEN_H_N:I VCC_IO:I VGND_IO:I
Xmpin_slow_q0 PD_I2C_H DRVLO_H_N int_slow VCC_IO sky130_fd_pr__pfet_g5v0d10v5
+ m=1 w=0.42 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpen_slow_q0 int_slow PDEN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=0.42 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpin_fast<1>_q0 PD_I2C_H DRVLO_H_N net62 VCC_IO sky130_fd_pr__pfet_g5v0d10v5
+ m=1 w=0.42 l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpin_fast<0>_q0 PD_I2C_H DRVLO_H_N net62 VCC_IO sky130_fd_pr__pfet_g5v0d10v5
+ m=1 w=0.42 l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpen_fast1_q0 net62 EN_FAST_N[1] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=0.42 l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI72<1> net53<0> EN_FAST_N[1] net42 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=3.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI72<0> net53<1> EN_FAST_N[0] net42 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=3.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI74<1> PD_H DRVLO_H_N net53<0> VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI74<0> PD_H DRVLO_H_N net53<1> VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI75 net039 PDEN_H_N net42 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=4.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI76 PD_H DRVLO_H_N net45 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=4.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI73 net42 I2C_MODE_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=3 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI101 net45 PDEN_H_N net039 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=4.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI94 PD_H I2C_MODE_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmnin_q0 PD_I2C_H DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2
+ w=3.0 l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnen_q0 PD_I2C_H PDEN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=3.0 l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI78 PD_H PDEN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI77 PD_H DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.6
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_pdpredrvr_strong_nr2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_pdpredrvr_strong_nr3 DRVLO_H_N EN_FAST_N[1]
+ EN_FAST_N[0] I2C_MODE_H PD_H PDEN_H_N VCC_IO VGND_IO
*.PININFO DRVLO_H_N:I EN_FAST_N[1]:I EN_FAST_N[0]:I I2C_MODE_H:I
*.PININFO PD_H:O PDEN_H_N:I VCC_IO:I VGND_IO:I
XI85 int1 I2C_MODE_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmpin_slow_q0 PD_H DRVLO_H_N int_slow VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=0.42 l=2.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpen_slow_q0 int_slow PDEN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=0.42 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpin_fast<1>_q0 PD_H DRVLO_H_N int_nor<1> VCC_IO sky130_fd_pr__pfet_g5v0d10v5
+ m=1 w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpin_fast<0>_q0 PD_H DRVLO_H_N int_nor<0> VCC_IO sky130_fd_pr__pfet_g5v0d10v5
+ m=1 w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmpen_fast<1>_q0 int_nor<1> EN_FAST_N[1] VCC_IO VCC_IO
+ sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xmpen_fast<0>_q0 int_nor<0> EN_FAST_N[0] VCC_IO VCC_IO
+ sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
XI90 PD_H DRVLO_H_N net43 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=2.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI56 net43 PDEN_H_N int1 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=2.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI87<1> PD_H DRVLO_H_N int2 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI87<0> PD_H DRVLO_H_N int2 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI86<1> int2 EN_FAST_N[1] int1 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI86<0> int2 EN_FAST_N[0] int1 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmnin_q0 PD_H DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=5 w=3.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmnen_q0 PD_H PDEN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_pdpredrvr_strong_nr3

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_pupredrvr_strong DRVHI_H PU_H_N[3] PU_H_N[2] PUEN_H
+ SLOW_H_N VCC_IO VGND_IO
*.PININFO DRVHI_H:I PU_H_N[3]:O PU_H_N[2]:O PUEN_H:I SLOW_H_N:I
*.PININFO VCC_IO:I VGND_IO:I
Xnd2b_q0 DRVHI_H en_fast_h_3<3> en_fast_h_3<2> en_fast_h_3<1> en_fast_h_3<0>
+ PU_H_N[3] PUEN_H VCC_IO VGND_IO sky130_fd_io__gpiov2_pupredrvr_strong_nd2
Xnd2a_q0 DRVHI_H net54 net54 net54 net54 PU_H_N[2] PUEN_H VCC_IO VGND_IO
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2
XI98 en_fast_h_3<0> en_fast_h_3<3> VGND_IO sky130_fd_io__tk_opti
XI97 en_fast_h_3<1> en_fast_h_3<3> VGND_IO sky130_fd_io__tk_opti
XI92 en_fast_h_3<3> nbias_out en_fast_h sky130_fd_io__tk_opto
XI96 en_fast_h_3<2> en_fast_h_3<3> VGND_IO sky130_fd_io__tk_opto
XI93 net54 nbias_out en_fast_h sky130_fd_io__tk_opto
Xinv_q0 en_fast_h_n en_fast_h VGND_IO VCC_IO sky130_fd_io__com_inv_x1_dnw
Xnbias_q0 DRVHI_H en_fast_h en_fast_h_n nbias_out PU_H_N[2] PUEN_H VCC_IO
+ VGND_IO sky130_fd_io__com_pupredrvr_nbias
Xnand_q0 PUEN_H SLOW_H_N en_fast_h_n VGND_IO VCC_IO sky130_fd_io__com_nand2_dnw
.ENDS sky130_fd_io__gpiov2_pupredrvr_strong

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_pupredrvr_strong_nd2 DRVHI_H EN_FAST[3] EN_FAST[2]
+ EN_FAST[1] EN_FAST[0] PU_H_N PUEN_H VCC_IO VGND_IO
*.PININFO DRVHI_H:I EN_FAST[3]:I EN_FAST[2]:I EN_FAST[1]:I
*.PININFO EN_FAST[0]:I PU_H_N:O PUEN_H:I VCC_IO:I VGND_IO:I
XE1 net24 PU_H_N sky130_fd_io__tk_em1s
Rrespu1 int_res net24 sky130_fd_pr__res_generic_po W=0.33 L=11 m=1
Rrespu2 PU_H_N int_res sky130_fd_pr__res_generic_po W=0.33 L=4 m=1
Xmnin_fast<3>_q0 net24 DRVHI_H int<3> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnin_fast<2>_q0 net24 DRVHI_H int<2> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnin_fast<1>_q0 net24 DRVHI_H int<1> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnin_fast<0>_q0 net24 DRVHI_H int<0> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnen_slow1_q0 n<2> PUEN_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=0.42 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnin_slow_q0 PU_H_N DRVHI_H n<2> VGND_IO sky130_fd_pr__nfet_g5v0d10v5 m=1
+ w=0.42 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xmnen_fast<3>_q0 int<3> EN_FAST[3] VGND_IO VGND_IO
+ sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xmnen_fast<2>_q0 int<2> EN_FAST[2] VGND_IO VGND_IO
+ sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xmnen_fast<1>_q0 int<1> EN_FAST[1] VGND_IO VGND_IO
+ sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xmnen_fast<0>_q0 int<0> EN_FAST[0] VGND_IO VGND_IO
+ sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.5 l=1.0 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xmpen_q0 PU_H_N PUEN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xmpin_q0 PU_H_N DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=3 w=5.0
+ l=0.6 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_pupredrvr_strong_nd2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__gpiov2_vcchib_in_buf IN_H MODE_VCCHIB_LV_N OUT OUT_N
+ VCCHIB VSSD
*.PININFO IN_H:I MODE_VCCHIB_LV_N:I OUT:O OUT_N:O VCCHIB:I VSSD:I
XI420 net57 in_b fbk VSSD sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI552 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI544 fbk IN_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI551 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI424 net81 in_b VSSD VSSD sky130_fd_pr__nfet_01v8 m=2 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI423 OUT_N net81 VSSD VSSD sky130_fd_pr__nfet_01v8 m=1 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI545 in_b IN_H fbk VSSD sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI487 OUT OUT_N VSSD VSSD sky130_fd_pr__nfet_01v8 m=3 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI541 net81 MODE_VCCHIB_LV_N VSSD VSSD sky130_fd_pr__nfet_01v8 m=2 w=1.0 l=0.25
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI549 net57 MODE_VCCHIB_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 m=1 w=5.0
+ l=0.25 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI436 net81 in_b net112 VCCHIB sky130_fd_pr__pfet_01v8 m=2 w=1.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI543 in_b IN_H net108 VCCHIB sky130_fd_pr__pfet_g5v0d10v5 m=2 w=5.0 l=0.8
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI429 OUT_N net81 VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 m=1 w=5.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI538 net112 MODE_VCCHIB_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 m=1 w=3.0
+ l=0.25 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI489 OUT OUT_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 m=1 w=5.0 l=0.25 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI547 net108 MODE_VCCHIB_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 m=3 w=5.0
+ l=0.25 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__gpiov2_vcchib_in_buf

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__hvsbt_inv_x1 IN OUT VGND VPWR
*.PININFO IN:I OUT:O VGND:I VPWR:I
XI1 OUT IN VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 OUT IN VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__hvsbt_inv_x1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__hvsbt_inv_x2 IN OUT VGND VPWR
*.PININFO IN:I OUT:O VGND:I VPWR:I
XI2 OUT IN VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__hvsbt_inv_x2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__hvsbt_inv_x4 IN OUT VGND VPWR
*.PININFO IN:I OUT:O VGND:I VPWR:I
XI1 OUT IN VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=8 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 OUT IN VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=4 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__hvsbt_inv_x4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__hvsbt_inv_x8 IN OUT VGND VPWR
*.PININFO IN:I OUT:O VGND:I VPWR:I
XI2 OUT IN VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=8 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=16 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__hvsbt_inv_x8

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__hvsbt_nand2 IN0 IN1 OUT VGND VPWR
*.PININFO IN0:I IN1:I OUT:O VGND:I VPWR:I
XI3 OUT IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI5 OUT IN1 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN1 net25 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 net25 IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__hvsbt_nand2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__hvsbt_nor IN0 IN1 OUT VGND VPWR
*.PININFO IN0:I IN1:I OUT:O VGND:I VPWR:I
XI3 net16 IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=2
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 OUT IN1 net16 VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=2
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 OUT IN1 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__hvsbt_nor

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__hvsbt_xor IN0 IN1 OUT VGND VPWR
*.PININFO IN0:I IN1:I OUT:O VGND:I VPWR:I
XI3 net29 IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI5 OUT net54 net45 VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI17 net70 IN1 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI18 net54 IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI13 net45 IN1 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 OUT net70 net29 VPWR sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN1 net58 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI16 net70 IN1 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 OUT net70 net62 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI15 net62 net54 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI14 net58 IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI19 net54 IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__hvsbt_xor

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__inv_1 A Y VGND VNB VPB VPWR
*.PININFO A:I Y:O VGND:I VNB:I VPB:I VPWR:I
XMIN1 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMIP1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__inv_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__nand2_1 A B Y VGND VNB VPB VPWR
*.PININFO A:I B:I Y:O VGND:I VNB:I VPB:I VPWR:I
XMP0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMP1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMN0 Y A sndA VNB sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMN1 sndA B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__nand2_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__nand2_2_enhpath IN0 IN1 OUT VGND VPWR
*.PININFO IN0:I IN1:I OUT:O VGND:I VPWR:I
XI3 OUT IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI5 OUT IN1 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=4 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN1 net25 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 net25 IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__nand2_2_enhpath

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__nor2_1 A B Y VGND VNB VPB VPWR
*.PININFO A:I B:I Y:O VGND:I VNB:I VPB:I VPWR:I
XMP0 VPWR A sndPA VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMP1 sndPA B Y VPB sky130_fd_pr__pfet_01v8_hvt m=1 w=1.12 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMN0 Y A VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMN1 Y B VGND VNB sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__nor2_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__nor2_4_enhpath IN0 IN1 OUT VGND VPWR
*.PININFO IN0:I IN1:I OUT:O VGND:I VPWR:I
XI3 net16 IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=16 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 OUT IN1 net16 VPWR sky130_fd_pr__pfet_g5v0d10v5 m=16 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=8 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 OUT IN1 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=8 w=0.7 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__nor2_4_enhpath

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__nor3_dnw IN0 IN1 IN2 OUT VGND VPWR
*.PININFO IN0:I IN1:I IN2:I OUT:O VGND:I VPWR:I
XI3 net43 IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 net39 IN1 net43 VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI16 OUT IN2 net39 VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 OUT IN1 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI18 OUT IN2 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__nor3_dnw

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__res250only_small PAD ROUT
*.PININFO PAD:B ROUT:B

* NOTE: Removed all but the primary resistor;  the other devices do not
* show up in the layout.
*
* RI175 net12 net16 sky130_fd_pr__res_generic_po W=2 L=10.07 m=1
* RI229 net16 ROUT sky130_fd_pr__res_generic_po W=2 L=0.17 m=1
* RI228 PAD net12 sky130_fd_pr__res_generic_po W=2 L=0.17 m=1
* RI237<1> net16 ROUT short
* RI237<2> net16 ROUT short
* RI234<1> PAD net12 short
* RI234<2> PAD net12 short
R0 PAD PAD sky130_fd_pr__res_generic_l1 w=0.27 l=0.005
R9 PAD PAD sky130_fd_pr__res_generic_l1 w=0.23 l=0.005
R5 PAD PAD sky130_fd_pr__res_generic_m1 w=2.01 l=0.01
R3 PAD PAD sky130_fd_pr__res_generic_po w=0.34 l=0.085
R7 PAD PAD sky130_fd_pr__res_generic_po w=0.3 l=0.085
R2 PAD ROUT sky130_fd_pr__res_generic_po w=2 l=10.07
R1 ROUT ROUT sky130_fd_pr__res_generic_l1 w=0.23 l=0.005
R10 ROUT ROUT sky130_fd_pr__res_generic_l1 w=0.27 l=0.005
R6 ROUT ROUT sky130_fd_pr__res_generic_m1 w=2.01 l=0.01
R4 ROUT ROUT sky130_fd_pr__res_generic_po w=0.34 l=0.085
R8 ROUT ROUT sky130_fd_pr__res_generic_po w=0.3 l=0.085

*RI175 PAD ROUT sky130_fd_pr__res_generic_po W=2 L=10.07 m=1
.ENDS sky130_fd_io__res250only_small

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__res75only_small PAD ROUT
*.PININFO PAD:B ROUT:B
RI175 PAD ROUT sky130_fd_pr__res_generic_po W=2 L=3.15 m=1
.ENDS sky130_fd_io__res75only_small

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

* Modified by Tim:  The resistors here are in an annular shape, and they overlap
* between cells such that the center of the resistor connects between the two
* devices.  To be correct, these two nets must come out as pins.

.SUBCKT sky130_fd_io__signal_5_sym_hv_local_5term GATE IN NBODY NWELLRING VGND net16
*.PININFO GATE:I IN:B NBODY:B NWELLRING:B VGND:B
XI1 IN GATE VGND NBODY sky130_fd_pr__esd_nfet_g5v0d10v5 m=1 w=5.4 l=0.6 mult=1
+ sa=0.0 sb=0.0 sd=0.0 topography=normal area=0.048 perim=0.94
* RI9 net18 NBODY short
* RI8 net16 NWELLRING short
RI9 net18 NBODY sky130_fd_pr__res_generic_m1 W=0.02 L=0.005
*RI8 net16 NWELLRING sky130_fd_pr__res_generic_m1 W=0.02 L=0.005
RI8 net16_ NWELLRING sky130_fd_pr__res_generic_m1 W=0.02 L=0.005
.ENDS sky130_fd_io__signal_5_sym_hv_local_5term

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__sio_hotswap_dly IN OUT OUT_N VCC_IO VGND
*.PININFO IN:I OUT:O OUT_N:O VCC_IO:I VGND:I
XI228 OUT_N a5 sky130_fd_io__tk_em1o
XI229 OUT_N a7 sky130_fd_io__tk_em1o
XI227 a6 OUT sky130_fd_io__tk_em1o
XI214 OUT_N a1 sky130_fd_io__tk_em1o
XI215 a2 OUT sky130_fd_io__tk_em1o
XEdly0 IN OUT sky130_fd_io__tk_em1o
XI217 OUT_N a3 sky130_fd_io__tk_em1s
XEdly2 a4 OUT sky130_fd_io__tk_em1s
XI196 a1 IN VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI204 a4 a3 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI199 a2 a1 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI198 a3 a2 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI232 a5 a4 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI231 a6 a5 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI230 a7 a6 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI197 a1 IN VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI202 a4 a3 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI201 a2 a1 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI200 a3 a2 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI235 a5 a4 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI234 a6 a5 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI233 a7 a6 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__sio_hotswap_dly

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__sio_hotswap_hys IN OUT VCC_IO VGND
*.PININFO IN:I OUT:O VCC_IO:I VGND:I
XI650 vcc_io_buf OUT int_n VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI649 int_n IN VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI648 OUT IN int_n VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=0.42 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI655 vgnd_buf VCC_IO VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI647 vgnd_buf OUT int_p VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI656 vcc_io_buf VGND VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI646 OUT IN int_p VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=2 w=1.5 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI645 int_p IN VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.5 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__sio_hotswap_hys

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__sio_hotswap_log_i2c_fix DISHS_H DISHS_H_N EN_H ENHS_H
+ ENHS_H_N ENHS_LAT_H_N EXITHS_H FORCEHI_H[1] OD_I_H_N VCC_IO VGND
*.PININFO DISHS_H:O DISHS_H_N:O EN_H:I ENHS_H:O ENHS_H_N:O
*.PININFO ENHS_LAT_H_N:I EXITHS_H:O FORCEHI_H[1]:I OD_I_H_N:I VCC_IO:I
*.PININFO VGND:I
XI664 net39 net46 DISHS_H VGND VGND VCC_IO VCC_IO sky130_fd_io__sio_hvsbt_nand2
XI663 net80 FORCEHI_H[1] net46 VGND VGND VCC_IO VCC_IO
+ sky130_fd_io__sio_hvsbt_nand2
XI662 OD_I_H_N EN_H net39 VGND VGND VCC_IO VCC_IO sky130_fd_io__sio_hvsbt_nand2
XI658 OD_I_H_N net80 VGND VGND VCC_IO VCC_IO sky130_fd_io__sio_hvsbt_inv_x1
XI666 ENHS_LAT_H_N net74 VGND VGND VCC_IO VCC_IO sky130_fd_io__sio_hvsbt_inv_x1
XI565 net74 ENHS_H_N VGND VGND VCC_IO VCC_IO sky130_fd_io__sio_hvsbt_inv_x1
XI667 DISHS_H DISHS_H_N VGND VGND VCC_IO VCC_IO sky130_fd_io__sio_hvsbt_inv_x1
XI637 ENHS_H_N ENHS_H VGND VGND VCC_IO VCC_IO sky130_fd_io__sio_hvsbt_inv_x1
XI553 net74 enhs_dly_h_n EXITHS_H VGND VGND VCC_IO VCC_IO
+ sky130_fd_io__sio_hvsbt_nor
XI521 net74 enhs_dly_h enhs_dly_h_n VCC_IO VGND sky130_fd_io__sio_hotswap_dly
.ENDS sky130_fd_io__sio_hotswap_log_i2c_fix

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__sio_hotswap_pghspd IN1 IN2 OUT VGND
*.PININFO IN1:I IN2:I OUT:O VGND:I
XEin2b VGND net25 sky130_fd_io__tk_em1o
XEoutb net38 OUT sky130_fd_io__tk_em1o
XEin1b VGND net27 sky130_fd_io__tk_em1o
XEin1a IN1 net27 sky130_fd_io__tk_em1s
XEouta net42 OUT sky130_fd_io__tk_em1s
XEin2a IN2 net25 sky130_fd_io__tk_em1s
XI481 net50 IN2 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI507 OUT IN1 net50 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI651 net42 net27 net34 VGND sky130_fd_pr__nfet_g5v0d10v5 m=6 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI654 net38 net27 net30 VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI652 net34 net25 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=6 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI653 net30 net25 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__sio_hotswap_pghspd

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__sio_hotswap_wpd E_N OUT VGND
*.PININFO E_N:I OUT:O VGND:I
XI198 npd<15> npd<16> sky130_fd_io__tk_em1o
XI209 VGND npd<14> sky130_fd_io__tk_em1o
XI196 npd<17> npd<18> sky130_fd_io__tk_em1o
XI197 npd<16> npd<17> sky130_fd_io__tk_em1o
XE20 npd<18> OUT sky130_fd_io__tk_em1o
XI208 npd<14> npd<15> sky130_fd_io__tk_em1o
Xnen17_q0 npd<17> E_N npd<16> VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xnen15_q0 npd<15> E_N npd<14> VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xnen14_q0 npd<14> E_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xnen16_q0 npd<16> E_N npd<15> VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xnen19_q0 OUT E_N npd<18> VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
Xnen18_q0 npd<18> E_N npd<17> VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=8.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__sio_hotswap_wpd

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__sio_hvsbt_inv_x1 IN OUT VGND VNB VPB VPWR
*.PININFO IN:I OUT:O VGND:I VNB:I VPB:I VPWR:I
XI2 OUT IN VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__sio_hvsbt_inv_x1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__sio_hvsbt_inv_x2 IN OUT VGND VNB VPB VPWR
*.PININFO IN:I OUT:O VGND:I VNB:I VPB:I VPWR:I
XI1 OUT IN VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=2 w=3.0 l=0.6 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 OUT IN VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=2 w=1.0 l=0.6 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__sio_hvsbt_inv_x2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__sio_hvsbt_inv_x4 IN OUT VGND VNB VPB VPWR
*.PININFO IN:I OUT:O VGND:I VNB:I VPB:I VPWR:I
XI2 OUT IN VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=4 w=1.0 l=0.6 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=4 w=3.0 l=0.6 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__sio_hvsbt_inv_x4

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__sio_hvsbt_nand2 IN0 IN1 OUT VGND VNB VPB VPWR
*.PININFO IN0:I IN1:I OUT:O VGND:I VNB:I VPB:I VPWR:I
XI3 OUT IN0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI5 OUT IN1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN1 net25 VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 net25 IN0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__sio_hvsbt_nand2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__sio_hvsbt_nor IN0 IN1 OUT VGND VNB VPB VPWR
*.PININFO IN0:I IN1:I OUT:O VGND:I VNB:I VPB:I VPWR:I
XI3 net17 IN0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI12 OUT IN1 net17 VPB sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI1 OUT IN0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 OUT IN1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.6 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__sio_hvsbt_nor

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__sio_tk_em1o A B
*.PININFO A:B B:B
RI1 A net11 short
RI2 B net7 short
.ENDS sky130_fd_io__sio_tk_em1o

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__sio_tk_em1s A B
*.PININFO A:B B:B
RI1 A net8 short
RI2 B net8 short
.ENDS sky130_fd_io__sio_tk_em1s

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__sio_tk_tie_r_out_esd A B
*.PININFO A:B B:B
Resd_r A B sky130_fd_pr__res_generic_po W=0.5 L=10.2 m=1
.ENDS sky130_fd_io__sio_tk_tie_r_out_esd

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__tk_em1o A B
*.PININFO A:B B:B
* RI1 A net11 short
* RI2 B net7 short
RI1 A net11 sky130_fd_pr__res_generic_m1 W=0.66 L=0.01
RI2 B net7 sky130_fd_pr__res_generic_m1 W=0.66 L=0.01
.ENDS sky130_fd_io__tk_em1o


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__tk_em1s A B
*.PININFO A:B B:B
* RI1 A net8 short
* RI2 B net8 short
RI1 A net8 sky130_fd_pr__res_generic_m1 W=0.66 L=0.01
RI2 B net8 sky130_fd_pr__res_generic_m1 W=0.66 L=0.01
.ENDS sky130_fd_io__tk_em1s


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__tk_em2o A B
*.PININFO A:B B:B
* RI1 A net11 short
* RI2 B net7 short
RI1 A net11 sky130_fd_pr__res_generic_m2 W=0.26 L=0.01
RI2 B net7 sky130_fd_pr__res_generic_m2 W=0.26 L=0.01
.ENDS sky130_fd_io__tk_em2o

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__tk_em2s A B
*.PININFO A:B B:B
* RI1 A net8 short
* RI2 B net8 short
RI1 A net8 sky130_fd_pr__res_generic_m2 W=0.26 L=0.01
RI2 B net8 sky130_fd_pr__res_generic_m2 W=0.26 L=0.01
.ENDS sky130_fd_io__tk_em2s

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__tk_opti OUT SPD SPU
*.PININFO OUT:B SPD:B SPU:B
Xe2_q0 SPD OUT sky130_fd_io__tk_em1o
Xe1_q0 OUT SPU sky130_fd_io__tk_em1s
.ENDS sky130_fd_io__tk_opti


* optiA is the same as opti, but uses tk_em2s, which is like tk_em1s
* but with a m2 short instead of a m1 short.

.SUBCKT sky130_fd_io__tk_optiA OUT SPD SPU
*.PININFO OUT:B SPD:B SPU:B
Xe2_q0 SPD OUT sky130_fd_io__tk_em1o
Xe1_q0 OUT SPU sky130_fd_io__tk_em2s
.ENDS sky130_fd_io__tk_optiA


* optiB is the same as opti, but uses tk_em2s, which is like tk_em1s
* but with a m2 short instead of a m1 short, and tk_em2o, which is
* like tk_em1o but with m2 shorts instead of m1 shorts.

.SUBCKT sky130_fd_io__tk_optiB OUT SPD SPU
*.PININFO OUT:B SPD:B SPU:B
Xe2_q0 SPD OUT sky130_fd_io__tk_em2o
Xe1_q0 OUT SPU sky130_fd_io__tk_em2s
.ENDS sky130_fd_io__tk_optiB


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__tk_opto OUT SPD SPU
*.PININFO OUT:B SPD:B SPU:B
Xe1_q0 SPU OUT sky130_fd_io__tk_em1o
Xe2_q0 OUT SPD sky130_fd_io__tk_em1s
.ENDS sky130_fd_io__tk_opto

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__tk_tie_r_out_esd A B
*.PININFO A:B B:B
Resd_r A B sky130_fd_pr__res_generic_po W=0.5 L=10.2 m=1
.ENDS sky130_fd_io__tk_tie_r_out_esd

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__top_amuxsplitv2 AMUXBUS_A_L AMUXBUS_A_R AMUXBUS_B_L
+ AMUXBUS_B_R ENABLE_VDDA_H HLD_VDDA_H_N SWITCH_AA_S0 SWITCH_AA_SL SWITCH_AA_SR
+ SWITCH_BB_S0 SWITCH_BB_SL SWITCH_BB_SR VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD
+ VSSIO VSSIO_Q VSWITCH
*.PININFO AMUXBUS_A_L:B AMUXBUS_A_R:B AMUXBUS_B_L:B AMUXBUS_B_R:B
*.PININFO ENABLE_VDDA_H:I HLD_VDDA_H_N:I SWITCH_AA_S0:I SWITCH_AA_SL:I
*.PININFO SWITCH_AA_SR:I SWITCH_BB_S0:I SWITCH_BB_SL:I SWITCH_BB_SR:I
*.PININFO VCCD:B VCCHIB:B VDDA:B VDDIO:B VDDIO_Q:B VSSA:B VSSD:B
*.PININFO VSSIO:B VSSIO_Q:B VSWITCH:B
xI22 VSSA VDDA sky130_fd_io__condiode
XI18 hold SWITCH_AA_S0 ng_vdda_aa_s0_h reset VCCD VDDA VSSA VSSD
+ sky130_fd_io__amuxsplitv2_switch_s0
XI348 hold SWITCH_BB_S0 ng_vdda_bb_s0_h reset VCCD VDDA VSSA VSSD
+ sky130_fd_io__amuxsplitv2_switch_s0
XI347 hold SWITCH_AA_SL ng_vswitch_aa_sl_h pg_vdda_aa_sl_h_n reset VCCD VDDA
+ VSSA VSSD VSWITCH sky130_fd_io__amuxsplitv2_switch_sl
XI24 hold SWITCH_AA_SR ng_vswitch_aa_sr_h pg_vdda_aa_sr_h_n reset VCCD VDDA VSSA
+ VSSD VSWITCH sky130_fd_io__amuxsplitv2_switch_sl
XI349 hold SWITCH_BB_SR ng_vswitch_bb_sr_h pg_vdda_bb_sr_h_n reset VCCD VDDA
+ VSSA VSSD VSWITCH sky130_fd_io__amuxsplitv2_switch_sl
XI350 hold SWITCH_BB_SL ng_vswitch_bb_sl_h pg_vdda_bb_sl_h_n reset VCCD VDDA
+ VSSA VSSD VSWITCH sky130_fd_io__amuxsplitv2_switch_sl
XI6 AMUXBUS_A_L AMUXBUS_A_R ng_vswitch_aa_sl_h ng_vswitch_aa_sr_h
+ ng_vdda_aa_s0_h pg_vdda_aa_sl_h_n pg_vdda_aa_sr_h_n VDDA VSSA
+ sky130_fd_io__amuxsplitv2_switch
XI8 AMUXBUS_B_L AMUXBUS_B_R ng_vswitch_bb_sl_h ng_vswitch_bb_sr_h
+ ng_vdda_bb_s0_h pg_vdda_bb_sl_h_n pg_vdda_bb_sr_h_n VDDA VSSA
+ sky130_fd_io__amuxsplitv2_switch
XI342 ENABLE_VDDA_H HLD_VDDA_H_N hold reset VDDA VSSA
+ sky130_fd_io__amuxsplitv2_delay
.ENDS sky130_fd_io__top_amuxsplitv2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__top_gpio_ovtv2 AMUXBUS_A AMUXBUS_B ANALOG_EN ANALOG_POL
+ ANALOG_SEL DM[2] DM[1] DM[0] ENABLE_H ENABLE_INP_H ENABLE_VDDA_H ENABLE_VDDIO
+ ENABLE_VSWITCH_H HLD_H_N HLD_OVR HYS_TRIM IB_MODE_SEL[1] IB_MODE_SEL[0] IN IN_H
+ INP_DIS OE_N OUT PAD PAD_A_ESD_0_H PAD_A_ESD_1_H PAD_A_NOESD_H SLEW_CTL[1]
+ SLEW_CTL[0] SLOW TIE_HI_ESD TIE_LO_ESD VCCD VCCHIB VDDA VDDIO VDDIO_Q VINREF
+ VSSA VSSD VSSIO VSSIO_Q VSWITCH VTRIP_SEL
*.PININFO AMUXBUS_A:B AMUXBUS_B:B ANALOG_EN:I ANALOG_POL:I
*.PININFO ANALOG_SEL:I DM[2]:I DM[1]:I DM[0]:I ENABLE_H:I
*.PININFO ENABLE_INP_H:I ENABLE_VDDA_H:I ENABLE_VDDIO:I
*.PININFO ENABLE_VSWITCH_H:I HLD_H_N:I HLD_OVR:I HYS_TRIM:I
*.PININFO IB_MODE_SEL[1]:I IB_MODE_SEL[0]:I IN:O IN_H:O INP_DIS:I
*.PININFO OE_N:I OUT:I PAD:B PAD_A_ESD_0_H:B PAD_A_ESD_1_H:B
*.PININFO PAD_A_NOESD_H:B SLEW_CTL[1]:I SLEW_CTL[0]:I SLOW:I
*.PININFO TIE_HI_ESD:O TIE_LO_ESD:O VCCD:B VCCHIB:B VDDA:B VDDIO:B
*.PININFO VDDIO_Q:B VINREF:I VSSA:B VSSD:B VSSIO:B VSSIO_Q:B VSWITCH:B
*.PININFO VTRIP_SEL:I
Xopath_q0 dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> hld_i_h_n
+ hld_i_ovr_h nga_pad_vpmp_h ngb_pad_vpmp_h od_i_h_n OE_N OUT PAD pd_csd_h pghs_h
+ pu_csd_h pug_h<6> pug_h<5> slew_ctl_h<1> slew_ctl_h<0> slew_ctl_h_n<1>
+ slew_ctl_h_n<0> SLOW TIE_HI_ESD TIE_LO_ESD VCCD VDDIO VDDIO_Q vpb_drvr VCCHIB
+ VSSA VSSD VSSIO VSSIO_Q sky130_fd_io__gpio_ovtv2_opath_i2c_fix_leak_fix
Xovt_amux_q0 AMUXBUS_A AMUXBUS_B ANALOG_EN ANALOG_POL ANALOG_SEL ENABLE_VDDA_H
+ ENABLE_VSWITCH_H hld_i_h_n nga_pad_vpmp_h ngb_pad_vpmp_h TIE_HI_ESD OUT PAD
+ pd_csd_h pghs_h pu_csd_h pug_h<6> pug_h<5> VCCD VDDA VDDIO VDDIO_Q vpb_drvr VSSA
+ VSSD VSSIO VSWITCH sky130_fd_io__gpio_ovtv2_amux_i2c_fix
Xctrl_q0 DM[2] DM[1] DM[0] dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0>
+ ENABLE_H ENABLE_INP_H HLD_H_N hld_i_h_n hld_i_ovr_h HLD_OVR HYS_TRIM hyst_trim_h
+ net164 IB_MODE_SEL[1] IB_MODE_SEL[0] ib_mode_sel_h<1> ib_mode_sel_h<0> net166<0>
+ net166<1> INP_DIS inp_dis_h_n od_i_h_n SLEW_CTL[1] SLEW_CTL[0] slew_ctl_h<1>
+ slew_ctl_h<0> slew_ctl_h_n<1> slew_ctl_h_n<0> VCCD VDDIO_Q VSSD VTRIP_SEL
+ vtrip_sel_h sky130_fd_io__gpio_ctlv2_i2c_fix
XI336 net193 PAD_A_ESD_1_H sky130_fd_io__res75only_small
XI335 PAD net193 sky130_fd_io__res75only_small
XI334 net189 PAD_A_ESD_0_H sky130_fd_io__res75only_small
Xresd4_q0 PAD net189 sky130_fd_io__res75only_small
Xipath_q0 dm_h_n<2> dm_h_n<1> dm_h_n<0> ENABLE_VDDIO hyst_trim_h
+ ib_mode_sel_h<1> ib_mode_sel_h<0> inp_dis_h_n IN IN_H PAD VCCHIB VDDIO_Q VINREF
+ VSSD vtrip_sel_h sky130_fd_io__gpio_ovtv2_ipath
RS0 PAD PAD_A_NOESD_H short
.ENDS sky130_fd_io__top_gpio_ovtv2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__top_gpiov2 AMUXBUS_A AMUXBUS_B ANALOG_EN ANALOG_POL
+ ANALOG_SEL DM[2] DM[1] DM[0] ENABLE_H ENABLE_INP_H ENABLE_VDDA_H ENABLE_VDDIO
+ ENABLE_VSWITCH_H HLD_H_N HLD_OVR IB_MODE_SEL IN IN_H INP_DIS OE_N OUT PAD
+ PAD_A_ESD_0_H PAD_A_ESD_1_H PAD_A_NOESD_H SLOW TIE_HI_ESD TIE_LO_ESD VCCD VCCHIB
+ VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH VTRIP_SEL
*.PININFO AMUXBUS_A:B AMUXBUS_B:B ANALOG_EN:I ANALOG_POL:I
*.PININFO ANALOG_SEL:I DM[2]:I DM[1]:I DM[0]:I ENABLE_H:I
*.PININFO ENABLE_INP_H:I ENABLE_VDDA_H:I ENABLE_VDDIO:I
*.PININFO ENABLE_VSWITCH_H:I HLD_H_N:I HLD_OVR:I IB_MODE_SEL:I IN:O
*.PININFO IN_H:O INP_DIS:I OE_N:I OUT:I PAD:B PAD_A_ESD_0_H:B
*.PININFO PAD_A_ESD_1_H:B PAD_A_NOESD_H:B SLOW:I TIE_HI_ESD:O
*.PININFO TIE_LO_ESD:O VCCD:B VCCHIB:B VDDA:B VDDIO:B VDDIO_Q:B VSSA:B
*.PININFO VSSD:B VSSIO:B VSSIO_Q:B VSWITCH:B VTRIP_SEL:I
Xamux_q0 AMUXBUS_A AMUXBUS_B ANALOG_EN ANALOG_POL ANALOG_SEL ENABLE_VDDA_H
+ ENABLE_VSWITCH_H hld_i_h hld_i_h_n OUT PAD VCCD VDDA VDDIO_Q VSSA VSSD VSSIO_Q
+ VSWITCH sky130_fd_io__gpiov2_amux
Xopath_q0 dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> hld_i_h_n
+ hld_i_ovr_h od_i_h OE_N OUT PAD SLOW TIE_HI_ESD TIE_LO_ESD VDDIO VSSD VSSIO VCCD
+ VCCHIB sky130_fd_io__gpiov2_opath
Xctrl_q0 DM[2] DM[1] DM[0] dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0>
+ ENABLE_H ENABLE_INP_H HLD_H_N hld_i_h hld_i_h_n hld_i_ovr_h HLD_OVR IB_MODE_SEL
+ ib_mode_sel_h ib_mode_sel_h_n INP_DIS inp_dis_h_n od_i_h VDDIO_Q VSSD VCCD
+ VTRIP_SEL vtrip_sel_h vtrip_sel_h_n sky130_fd_io__gpiov2_ctl
Xipath_q0 dm_h_n<2> dm_h_n<1> dm_h_n<0> ENABLE_VDDIO ib_mode_sel_h
+ ib_mode_sel_h_n inp_dis_h_n IN IN_H PAD VCCHIB VDDIO_Q VSSD vtrip_sel_h_n
+ sky130_fd_io__gpiov2_ipath
Xresd3_q0 PAD_A_ESD_1_H net210 sky130_fd_io__res75only_small
Xresd1_q0 net204 PAD sky130_fd_io__res75only_small
Xresd4_q0 net210 PAD sky130_fd_io__res75only_small
Xresd2_q0 PAD_A_ESD_0_H net204 sky130_fd_io__res75only_small
* RS0<2> PAD PAD_A_NOESD_H short
* RS0<1> PAD PAD_A_NOESD_H short
* RS0<0> PAD PAD_A_NOESD_H short
RS0<2> PAD PAD_A_NOESD_H sky130_fd_pr__res_generic_m4 W=12.35 L=0.035
RS0<1> PAD PAD_A_NOESD_H sky130_fd_pr__res_generic_m3 W=1.07 L=0.035
RS0<0> PAD PAD_A_NOESD_H sky130_fd_pr__res_generic_m3 W=12.37 L=0.035
.ENDS sky130_fd_io__top_gpiov2


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__top_ground_hvc_wpad AMUXBUS_A AMUXBUS_B DRN_HVC G_CORE
+ G_PAD OGC_HVC PADISOL PADISOR SRC_BDY_HVC VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA
+ VSSD VSSIO VSSIO_Q VSWITCH
*.PININFO AMUXBUS_A:B AMUXBUS_B:B DRN_HVC:B G_CORE:B G_PAD:B OGC_HVC:B
*.PININFO PADISOL:B PADISOR:B SRC_BDY_HVC:B VCCD:B VCCHIB:B VDDA:B VDDIO:B
*.PININFO VDDIO_L:B VSSA:B VSSD:B VSSIO:B VSSIO_Q:B VSWITCH:B
xI39 SRC_BDY_HVC VDDIO sky130_fd_io__condiode
Xcxtor2_q0 DRN_HVC g_nclamp SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5
+ m=22 w=10.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xnc2_q0 SRC_BDY_HVC g_pdpre SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5
+ m=5 w=5.0 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xnc1_q0 SRC_BDY_HVC g_pdpre SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5
+ m=15 w=5.0 l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xpre_n1_q0 g_nclamp g_pdpre SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5
+ m=15 w=7.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xclamp_xtor_q0 DRN_HVC g_nclamp SRC_BDY_HVC SRC_BDY_HVC
+ sky130_fd_pr__nfet_g5v0d10v5 m=120 w=20.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Rrc_res g_pdpre net94 sky130_fd_pr__res_generic_po W=0.33 L=470 m=1
RI38 net90 DRN_HVC sky130_fd_pr__res_generic_po W=0.33 L=700 m=1
RI37 net94 net90 sky130_fd_pr__res_generic_po W=0.33 L=1550 m=1
Xpre_p1_q0 g_nclamp g_pdpre DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 m=50
+ w=7.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
RI13 G_PAD G_CORE sky130_fd_pr__res_generic_m5 w=2.5385e+08u l=100000u
RIL G_CORE PADISOL sky130_fd_pr__res_generic_m3 w=11.825 l=0.01
RIR G_CORE PADISOR sky130_fd_pr__res_generic_m3 w=11.825 l=0.01
.ENDS sky130_fd_io__top_ground_hvc_wpad

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__top_hvclamp_wopadv2 DRN_HVC OGC_HVC SRC_BDY_HVC VSSD
*.PININFO DRN_HVC:B OGC_HVC:B SRC_BDY_HVC:B VSSD:B
xI39 SRC_BDY_HVC OGC_HVC sky130_fd_io__condiode
Xpre_p1_q0 g_nclamp g_pdpre DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 m=50
+ w=7.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Rrc_res g_pdpre net41 sky130_fd_pr__res_generic_po W=0.33 L=470 m=1
RI38 net37 DRN_HVC sky130_fd_pr__res_generic_po W=0.33 L=700 m=1
RI37 net41 net37 sky130_fd_pr__res_generic_po W=0.33 L=1550 m=1
Xclamp_xtor_q0 DRN_HVC g_nclamp SRC_BDY_HVC SRC_BDY_HVC
+ sky130_fd_pr__nfet_g5v0d10v5 m=120 w=20.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xpre_n1_q0 g_nclamp g_pdpre SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5
+ m=15 w=7.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xnc1_q0 SRC_BDY_HVC g_pdpre SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5
+ m=15 w=5.0 l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xnc2_q0 SRC_BDY_HVC g_pdpre SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5
+ m=5 w=5.0 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xcxtor2_q0 DRN_HVC g_nclamp SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5
+ m=22 w=10.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
.ENDS sky130_fd_io__top_hvclamp_wopadv2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__top_power_hvc_wpadv2 AMUXBUS_A AMUXBUS_B DRN_HVC OGC_HVC
+ PADISOL PADISOR P_CORE P_PAD SRC_BDY_HVC VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA
+ VSSD VSSIO VSSIO_Q VSWITCH
*.PININFO AMUXBUS_A:B AMUXBUS_B:B DRN_HVC:B OGC_HVC:B PADISOL:B PADISOR:B
*.PININFO P_CORE:B P_PAD:B SRC_BDY_HVC:B VCCD:B VCCHIB:B VDDA:B VDDIO:B
*.PINFNFO VDDIO_Q:B VSSA:B VSSD:B VSSIO:B VSSIO_Q:B VSWITCH:B
xI39 SRC_BDY_HVC VDDIO sky130_fd_io__condiode
Xpre_p1_q0 g_nclamp g_pdpre DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 m=50
+ w=7.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Rrc_res g_pdpre net67 sky130_fd_pr__res_generic_po W=0.33 L=470 m=1
RI38 net63 DRN_HVC sky130_fd_pr__res_generic_po W=0.33 L=700 m=1
RI37 net67 net63 sky130_fd_pr__res_generic_po W=0.33 L=1550 m=1
Xclamp_xtor_q0 DRN_HVC g_nclamp SRC_BDY_HVC SRC_BDY_HVC
+ sky130_fd_pr__nfet_g5v0d10v5 m=120 w=20.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xpre_n1_q0 g_nclamp g_pdpre SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5
+ m=15 w=7.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xnc1_q0 SRC_BDY_HVC g_pdpre SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5
+ m=15 w=5.0 l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xnc2_q0 SRC_BDY_HVC g_pdpre SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5
+ m=5 w=5.0 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xcxtor2_q0 DRN_HVC g_nclamp SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5
+ m=22 w=10.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
RI13 P_PAD P_CORE sky130_fd_pr__res_generic_m5 w=2.5385e+08u l=100000u
RIL P_CORE PADISOL sky130_fd_pr__res_generic_m3 w=11.825 l=0.01
RIR P_CORE PADISOR sky130_fd_pr__res_generic_m3 w=11.825 l=0.01
.ENDS sky130_fd_io__top_power_hvc_wpadv2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__top_vrefcapv2 AMUXBUS_A AMUXBUS_B CNEG CPOS VCCD VCCHIB
+ VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH
*.PININFO AMUXBUS_A:B AMUXBUS_B:B CNEG:B CPOS:B VCCD:B VCCHIB:B VDDA:B
*.PININFO VDDIO:B VDDIO_Q:B VSSA:B VSSD:B VSSIO:B VSSIO_Q:B VSWITCH:B
xI271 CNEG VDDIO_Q sky130_fd_io__condiode
XI334 CNEG CPOS CNEG CNEG sky130_fd_pr__nfet_05v0_nvt m=180 w=10.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__top_vrefcapv2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

* Modified by Tim:  Split power and ground nets on XI364<1:0> fixed

.SUBCKT sky130_fd_io__top_xres4v2 AMUXBUS_A AMUXBUS_B DISABLE_PULLUP_H
+ EN_VDDIO_SIG_H ENABLE_H ENABLE_VDDIO FILT_IN_H INP_SEL_H PAD PAD_A_ESD_H
+ PULLUP_H TIE_HI_ESD TIE_LO_ESD TIE_WEAK_HI_H VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA
+ VSSD VSSIO VSSIO_Q VSWITCH XRES_H_N
*.PININFO AMUXBUS_A:B AMUXBUS_B:B DISABLE_PULLUP_H:I EN_VDDIO_SIG_H:I
*.PININFO ENABLE_H:I ENABLE_VDDIO:I FILT_IN_H:I INP_SEL_H:I PAD:B
*.PININFO PAD_A_ESD_H:B PULLUP_H:B TIE_HI_ESD:O TIE_LO_ESD:O
*.PININFO TIE_WEAK_HI_H:B VCCD:I VCCHIB:I VDDA:I VDDIO:I VDDIO_Q:I
*.PININFO VSSA:I VSSD:I VSSIO:I VSSIO_Q:I VSWITCH:I XRES_H_N:O
XI326 VSSIO TIE_LO_ESD sky130_fd_io__tk_tie_r_out_esd
XI49 VDDIO TIE_HI_ESD sky130_fd_io__tk_tie_r_out_esd
Xgpio_inbuf_q0 ENABLE_H ENABLE_VDDIO net79 net83 in_h VCCHIB VDDIO_Q VSSD
+ EN_VDDIO_SIG_H en_vddio_sig_h_n sky130_fd_io__xres4v2_in_buf
Xxresesd_q0 in_h net86 PAD VDDIO VSSD VSSIO sky130_fd_io__xres_esd
Xweakpullup_q0 TIE_WEAK_HI_H VDDIO VSSD sky130_fd_io__xres_wpu
Xesd_res_q0 PAD PAD_A_ESD_H sky130_fd_io__res250only_small
XI335 net97 PULLUP_H VSSD sky130_fd_io__com_xres_weak_pu
XI363 INP_SEL_H inp_sel_h_n VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x2
XI334 net103 net107 VSSD VDDIO sky130_fd_io__hvsbt_inv_x2
XI333 DISABLE_PULLUP_H net103 VSSD VDDIO sky130_fd_io__hvsbt_inv_x2
XI374 EN_VDDIO_SIG_H en_vddio_sig_h_n VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x2
XI368 net124 out_rcfilt_h VDDIO_Q VSSD sky130_fd_io__xres_rcfilter_lpf
XI367 out_rcfilt_h out_hysbuf_h VDDIO_Q VSSD sky130_fd_io__xres_inv_hys
XI365 out_hysbuf_h out_h_n VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x1
XI364<1> out_h_n XRES_H_N VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x4
XI364<0> out_h_n XRES_H_N VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x4
XI361 net124 inp_sel_h_n FILT_IN_H VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=3.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI358 net124 INP_SEL_H net79 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI332 net97 net107 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=4 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI360 net124 INP_SEL_H FILT_IN_H VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI357 net124 inp_sel_h_n net79 VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__top_xres4v2

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__xor2_1 A B X VGND VPWR
*.PININFO A:I B:I X:O VGND:I VPWR:I
XMNnor0 inor A VGND VGND sky130_fd_pr__nfet_01v8 m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMNnor1 inor B VGND VGND sky130_fd_pr__nfet_01v8 m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMNaoi10 VGND A sndNA VGND sky130_fd_pr__nfet_01v8 m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMNaoi11 sndNA B X VGND sky130_fd_pr__nfet_01v8 m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMNaoi20 X inor VGND VGND sky130_fd_pr__nfet_01v8 m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMPnor0 VPWR A sndPA VPWR sky130_fd_pr__pfet_01v8_hvt m=1 w=1.26 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMPnor1 sndPA B inor VPWR sky130_fd_pr__pfet_01v8_hvt m=1 w=1.26 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMPaoi10 pmid A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt m=1 w=1.26 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMPaoi11 pmid B VPWR VPWR sky130_fd_pr__pfet_01v8_hvt m=1 w=1.26 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XMPaoi20 X inor pmid VPWR sky130_fd_pr__pfet_01v8_hvt m=1 w=1.26 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__xor2_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__xres4v2_in_buf ENABLE_HV ENABLE_VDDIO_LV IN_H IN_H_N PAD
+ VCCHIB VDDIO VGND VNORMAL VNORMAL_B
*.PININFO ENABLE_HV:I ENABLE_VDDIO_LV:I IN_H:O IN_H_N:O PAD:I VCCHIB:I
*.PININFO VDDIO:I VGND:I VNORMAL:I VNORMAL_B:I
XI165 ENABLE_VDDIO_LV enable_vddio_lv_n VGND VGND VCCHIB VCCHIB
+ sky130_fd_io__inv_1
XI61 net106 mode_vcchib VGND VDDIO sky130_fd_io__hvsbt_inv_x1
XI35 VNORMAL_B ENABLE_HV net106 VGND VDDIO sky130_fd_io__hvsbt_nand2
XI132 net207 net110 VGND sky130_fd_pr__res_generic_nd__hv W=0.29 L=1077.19 m=1
RI159 net235 net108 sky130_fd_pr__res_generic_po W=0.4 L=713.695 m=1
XI8 net193 pad1 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI86 pad1 pad_inv VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI85 pad_inv PAD net140 VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI114 net152 pad_inv net140 VGND sky130_fd_pr__nfet_g5v0d10v5 m=4 w=5.0 l=0.8
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI145 enable_hv_b ENABLE_HV VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI251 IN_H IN_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=3 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI83 net140 PAD VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0 l=0.8 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI7 fbk pad_inv VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=2 w=5.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI213 IN_H_N fbk VGND VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI152 VGND VGND VGND VGND sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI113 net124 PAD net152 VGND sky130_fd_pr__nfet_05v0_nvt m=1 w=1.0 l=0.9 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI154 net120 mode_vcchib net206 VGND sky130_fd_pr__nfet_05v0_nvt m=1 w=1.0 l=0.9
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI151 net116 mode_vcchib vcchib_int VGND sky130_fd_pr__nfet_05v0_nvt m=1 w=10.0
+ l=0.9 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI150 net112 pad_inv net140 VGND sky130_fd_pr__nfet_g5v0d10v5 m=1 w=5.0 l=0.8
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI116 pad1 pad_inv net235 VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI143 net124 VNORMAL VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI156 net116 enable_vddio_lv_n VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI252 IN_H IN_H_N VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=3 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI107 net108 mode_vcchib VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI146 enable_hv_b ENABLE_HV VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI88 pad_inv PAD vcchib_int vcchib_int sky130_fd_pr__pfet_g5v0d10v5 m=1 w=1.0
+ l=0.8 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI89 pad_inv PAD net207 VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI90 pad1 pad_inv net206 net206 sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI133 net110 mode_vcchib VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0
+ l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI2 net193 fbk VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI219 fbk net193 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI14 IN_H_N fbk VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI158 net120 enable_vddio_lv_n VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 m=1
+ w=5.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI139 net207 VNORMAL_B net110 VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI136 net112 VNORMAL_B VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI153 vcchib_int vcchib_int vcchib_int vcchib_int sky130_fd_pr__pfet_g5v0d10v5
+ m=1 w=1.0 l=0.8 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI160 net235 VNORMAL_B net108 VDDIO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=5.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__xres4v2_in_buf

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__xres_esd OUT_H OUT_VT PAD VDDIO VSSD VSSIO
*.PININFO OUT_H:B OUT_VT:B PAD:B VDDIO:B VSSD:B VSSIO:B
Xesd_q0 PAD OUT_H OUT_VT VDDIO VSSD VSSD sky130_fd_io__gpio_buf_localesd
Xpddrvr_strong_q0 tie_lo_esd tie_lo_esd PAD tie_lo_esd tie_lo_esd tie_lo_esd
+ VDDIO VSSIO VSSIO sky130_fd_io__gpio_pddrvr_strong
Xpudrvr_strong_q0 PAD tie_hi_esd tie_hi_esd tie_hi_esd VDDIO VSSD
+ sky130_fd_io__gpio_pudrvr_strong
xI271 VSSIO VDDIO sky130_fd_io__condiode
.ENDS sky130_fd_io__xres_esd

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__xres_inv_hys IN_H OUT_H VCC_IO VSSD
*.PININFO IN_H:I OUT_H:O VCC_IO:I VSSD:I
XI7 pmid1 IN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI8 out_h_n IN_H pmid1 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI9 OUT_H out_h_n VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=3.0 l=0.5
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI10 pmid1 OUT_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 m=1 w=0.42 l=1.0
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI4 out_h_n IN_H nmid1 VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI5 nmid1 IN_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI6 OUT_H out_h_n VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=1.0 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI11 nmid1 OUT_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 m=1 w=0.42 l=1.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__xres_inv_hys

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__xres_rcfilter_lpf IN OUT VCC_IO VSSD
*.PININFO IN:I OUT:O VCC_IO:B VSSD:B
Xe5_q0 net65 net40 sky130_fd_io__xres_tk_emlo
Xe1_q0 net135 net67 sky130_fd_io__xres_tk_emlo
Xe4_q0 net43 net65 sky130_fd_io__xres_tk_emlo
XI200 net59 OUT sky130_fd_io__xres_tk_emlo
XI199 net62 OUT sky130_fd_io__xres_tk_emlo
XI198 VSSD net59 sky130_fd_io__xres_tk_emlo
XI197 VSSD net57 sky130_fd_io__xres_tk_emlo
XI194 net57 OUT sky130_fd_io__xres_tk_emlo
XI193 net45 OUT sky130_fd_io__xres_tk_emlo
XI191 net42 OUT sky130_fd_io__xres_tk_emlo
XI190 net40 OUT sky130_fd_io__xres_tk_emlo
XI187 VSSD OUT sky130_fd_io__xres_tk_emlo
XI186 VSSD net45 sky130_fd_io__xres_tk_emlo
Xe2_q0 net67 net43 sky130_fd_io__xres_tk_emlo
XI183 net42 VSSD sky130_fd_io__xres_tk_emlo
XI181 net40 VSSD sky130_fd_io__xres_tk_emlo
XI202 VSSD sky130_fd_io__xres_tk_emlc
XI201 VSSD sky130_fd_io__xres_tk_emlc
XI192 OUT sky130_fd_io__xres_tk_emlc
XI189 VSSD sky130_fd_io__xres_tk_emlc
XI188 VSSD sky130_fd_io__xres_tk_emlc
XI180 net40 sky130_fd_io__xres_tk_emlc
XI182 net42 sky130_fd_io__xres_tk_emlc
Xe3_q0 net43 sky130_fd_io__xres_tk_emlc
XI172 IN net135 VSSD VSSD VCC_IO sky130_fd_io__xres_rcfilter_lpf_rcunit
XI184 VSSD net57 VSSD VSSD VCC_IO sky130_fd_io__xres_rcfilter_lpf_rcunit
XI185 VSSD net45 VSSD VSSD VCC_IO sky130_fd_io__xres_rcfilter_lpf_rcunit
XI196 VSSD net62 VSSD VSSD VCC_IO sky130_fd_io__xres_rcfilter_lpf_rcunit
XI195 VSSD net59 VSSD VSSD VCC_IO sky130_fd_io__xres_rcfilter_lpf_rcunit
XI179 net43 net65 VSSD VSSD VCC_IO sky130_fd_io__xres_rcfilter_lpf_rcunit
XI178 net65 net40 VSSD VSSD VCC_IO sky130_fd_io__xres_rcfilter_lpf_rcunit
XI177 net40 net42 VSSD VSSD VCC_IO sky130_fd_io__xres_rcfilter_lpf_rcunit
XI176 net42 OUT VSSD VSSD VCC_IO sky130_fd_io__xres_rcfilter_lpf_rcunit
XI175 net67 net43 VSSD VSSD VCC_IO sky130_fd_io__xres_rcfilter_lpf_rcunit
XI174 net43 net43 VSSD VSSD VCC_IO sky130_fd_io__xres_rcfilter_lpf_rcunit
XI173 net135 net67 VSSD VSSD VCC_IO sky130_fd_io__xres_rcfilter_lpf_rcunit
.ENDS sky130_fd_io__xres_rcfilter_lpf

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__xres_rcfilter_lpf_rcunit IN OUT VGND VNB VPWR
*.PININFO IN:I OUT:O VGND:B VNB:B VPWR:B
Xr1b_q0 net14 OUT VNB sky130_fd_io__xres_rcfilter_lpf_res_sub
Xr1a_q0 IN net14 VNB sky130_fd_io__xres_rcfilter_lpf_res_sub
XI242 VGND OUT VGND VNB sky130_fd_pr__nfet_g5v0d10v5 m=1 w=7.0 l=4.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
XI244 VPWR OUT VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 m=1 w=7.0 l=4.0 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_io__xres_rcfilter_lpf_rcunit

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

* Modified by Tim:  Added 3rd terminal to sky130_fd_pr__res_generic_nd devices

.SUBCKT sky130_fd_io__xres_rcfilter_lpf_res_sub IN OUT VGND
*.PININFO IN:I OUT:O VGND:B
Xe1_q0 IN sky130_fd_io__xres_tk_emlc
Xe2_q0 OUT net30 sky130_fd_io__xres_tk_emlo
Xropti OUT net30 VGND sky130_fd_pr__res_generic_nd W=0.5 L=14 m=1
Xr1 net30 IN VGND sky130_fd_pr__res_generic_nd W=0.5 L=47 m=1
Xropto IN IN VGND sky130_fd_pr__res_generic_nd W=0.5 L=14 m=1
.ENDS sky130_fd_io__xres_rcfilter_lpf_res_sub

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__xres_tk_emlc A
*.PININFO A:B
* RI2 A net7 short
* RI1 A net2 short
RI2 A net7 sky130_fd_pr__res_generic_m1 W=0.66 L=0.01
RI1 A net2 sky130_fd_pr__res_generic_m1 W=0.66 L=0.01
.ENDS sky130_fd_io__xres_tk_emlc

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__xres_tk_emlo A B
*.PININFO A:B B:B
* RI2 B net8 short
* RI1 A net3 short
RI2 B net8 sky130_fd_pr__res_generic_m1 W=0.66 L=0.01
RI1 A net3 sky130_fd_pr__res_generic_m1 W=0.66 L=0.01
.ENDS sky130_fd_io__xres_tk_emlo

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__xres_wpu PAD VDDIO VSSD
*.PININFO PAD:B VDDIO:B VSSD:B
Xesdr_q0 PAD net15 sky130_fd_io__res250only_small
X5kres_q0 VDDIO net15 VSSD sky130_fd_io__com_res_weak
.ENDS sky130_fd_io__xres_wpu

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__top_ground_lvc_wpad AMUXBUS_A AMUXBUS_B BDY2_B2B DRN_LVC1
+ DRN_LVC2 G_CORE G_PAD OGC_LVC PADISOL PADISOR SRC_BDY_LVC1 SRC_BDY_LVC2 VCCD
+ VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH
*.PININFO AMUXBUS_A:B AMUXBUS_B:B BDY2_B2B:B DRN_LVC1:B DRN_LVC2:B
*.PININFO G_CORE:B G_PAD:B OGC_LVC:B PADISOL:B PADISOR:B SRC_BDY_LVC1:B
*.PININFO SRC_BDY_LVC2:B VCCD:B VCCHIB:B VDDA:B VDDIO:B VDDIO_Q:B VSSA:B
*.PININFO VSSD:B VSSIO:B VSSIO_Q:B VSWITCH:B
Xesd_q0 BDY2_B2B SRC_BDY_LVC1 VSSD sky130_fd_io__gnd2gnd_120x2_lv_isosub
xI54 SRC_BDY_LVC2 VDDIO sky130_fd_io__condiode
xI50 SRC_BDY_LVC1 VDDIO sky130_fd_io__condiode
RI21 G_PAD G_CORE sky130_fd_pr__res_generic_m5 w=2.5385e+08u l=100000u
RIL G_CORE PADISOL sky130_fd_pr__res_generic_m3 w=11.825 l=0.01
RIR G_CORE PADISOR sky130_fd_pr__res_generic_m3 w=11.825 l=0.01
Xpre_p1_q0 g_nclamp_lvc1 g_pdpre_lvc1 DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8
+ m=20 w=7.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI40 g_nclamp_lvc2 g_pdpre_lvc2 DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 m=20
+ w=7.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xclamp_xtor_q0 DRN_LVC1 g_nclamp_lvc1 SRC_BDY_LVC1 SRC_BDY_LVC1
+ sky130_fd_pr__nfet_01v8 m=166 w=7.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
XI42 DRN_LVC2 g_nclamp_lvc2 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8
+ m=152 w=7.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI61 DRN_LVC2 g_nclamp_lvc2 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8
+ m=38 w=5.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI62 DRN_LVC1 g_nclamp_lvc1 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8
+ m=20 w=5.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xncap_q0 SRC_BDY_LVC1 g_pdpre_lvc1 SRC_BDY_LVC1 SRC_BDY_LVC1
+ sky130_fd_pr__nfet_01v8 m=15 w=7.0 l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xpre_n1_q0 g_nclamp_lvc1 g_pdpre_lvc1 SRC_BDY_LVC1 SRC_BDY_LVC1
+ sky130_fd_pr__nfet_01v8 m=3 w=7.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
XI43 g_nclamp_lvc2 g_pdpre_lvc2 SRC_BDY_LVC2 SRC_BDY_LVC2
+ sky130_fd_pr__nfet_01v8 m=2 w=7.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
XI58 SRC_BDY_LVC2 g_pdpre_lvc2 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8
+ m=6 w=5.0 l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI60 SRC_BDY_LVC2 g_pdpre_lvc2 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8
+ m=1 w=5.0 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI59 SRC_BDY_LVC2 g_pdpre_lvc2 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8
+ m=10 w=7.0 l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Rrc_res g_pdpre_lvc1 DRN_LVC1 sky130_fd_pr__res_generic_po W=0.33 L=1950 m=1
RI44 DRN_LVC2 net161 sky130_fd_pr__res_generic_po W=0.33 L=900 m=1
RI47 net161 net155 sky130_fd_pr__res_generic_po W=0.33 L=300 m=1
RI46 g_pdpre_lvc2 net157 sky130_fd_pr__res_generic_po W=0.33 L=200 m=1
RI45 net157 net155 sky130_fd_pr__res_generic_po W=0.33 L=720 m=1
.ENDS sky130_fd_io__top_ground_lvc_wpad

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_io__top_power_lvc_wpad AMUXBUS_A AMUXBUS_B BDY2_B2B DRN_LVC1
+ DRN_LVC2 OGC_LVC PADISOL PADISOR P_CORE P_PAD SRC_BDY_LVC1 SRC_BDY_LVC2 VCCD
+ VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH
*.PININFO AMUXBUS_A:B AMUXBUS_B:B BDY2_B2B:B DRN_LVC1:B DRN_LVC2:B
*.PININFO OGC_LVC:B PADISOL:B PADISOR:B P_CORE:B P_PAD:B SRC_BDY_LVC1:B
*.PININFO SRC_BDY_LVC2:B VCCD:B VCCHIB:B VDDA:B VDDIO:B VDDIO_Q:B
*.PININFO VSSA:B VSSD:B VSSIO:B VSSIO_Q:B VSWITCH:B
Xesd_q0 BDY2_B2B SRC_BDY_LVC1 VSSD sky130_fd_io__gnd2gnd_120x2_lv_isosub
xI54 SRC_BDY_LVC2 VDDIO sky130_fd_io__condiode
xI50 SRC_BDY_LVC1 VDDIO sky130_fd_io__condiode
RI21 P_PAD P_CORE sky130_fd_pr__res_generic_m5 w=2.5385e+08u l=100000u
RIL P_CORE PADISOL sky130_fd_pr__res_generic_m3 w=11.825 l=0.01
RIR P_CORE PADISOR sky130_fd_pr__res_generic_m3 w=11.825 l=0.01
Xpre_p1_q0 g_nclamp_lvc1 g_pdpre_lvc1 DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8
+ m=20 w=7.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI40 g_nclamp_lvc2 g_pdpre_lvc2 DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 m=20
+ w=7.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xclamp_xtor_q0 DRN_LVC1 g_nclamp_lvc1 SRC_BDY_LVC1 SRC_BDY_LVC1
+ sky130_fd_pr__nfet_01v8 m=166 w=7.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
XI42 DRN_LVC2 g_nclamp_lvc2 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8
+ m=152 w=7.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI61 DRN_LVC2 g_nclamp_lvc2 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8
+ m=38 w=5.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI62 DRN_LVC1 g_nclamp_lvc1 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8
+ m=20 w=5.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Xncap_q0 SRC_BDY_LVC1 g_pdpre_lvc1 SRC_BDY_LVC1 SRC_BDY_LVC1
+ sky130_fd_pr__nfet_01v8 m=15 w=7.0 l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
Xpre_n1_q0 g_nclamp_lvc1 g_pdpre_lvc1 SRC_BDY_LVC1 SRC_BDY_LVC1
+ sky130_fd_pr__nfet_01v8 m=3 w=7.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
XI43 g_nclamp_lvc2 g_pdpre_lvc2 SRC_BDY_LVC2 SRC_BDY_LVC2
+ sky130_fd_pr__nfet_01v8 m=2 w=7.0 l=0.18 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
XI58 SRC_BDY_LVC2 g_pdpre_lvc2 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8
+ m=6 w=5.0 l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI60 SRC_BDY_LVC2 g_pdpre_lvc2 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8
+ m=1 w=5.0 l=4.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
XI59 SRC_BDY_LVC2 g_pdpre_lvc2 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8
+ m=10 w=7.0 l=8.0 mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
Rrc_res g_pdpre_lvc1 DRN_LVC1 sky130_fd_pr__res_generic_po W=0.33 L=1950 m=1
RI44 DRN_LVC2 net161 sky130_fd_pr__res_generic_po W=0.33 L=900 m=1
RI47 net161 net155 sky130_fd_pr__res_generic_po W=0.33 L=300 m=1
RI46 g_pdpre_lvc2 net157 sky130_fd_pr__res_generic_po W=0.33 L=200 m=1
RI45 net157 net155 sky130_fd_pr__res_generic_po W=0.33 L=720 m=1
.ENDS sky130_fd_io__top_power_lvc_wpad
